************************************************************************
* auCdl Netlist:
* 
* Library Name:  VLSI
* Top Cell Name: DFFTG
* View Name:     schematic
* Netlisted on:  Nov 16 16:50:23 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: VLSI
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG A B EN ENbar VDD VSS
*.PININFO EN:I ENbar:I A:B B:B VDD:B VSS:B
MM1 A ENbar B VDD p_18 W=1u L=180.00n m=1
MM0 A EN B VSS n_18 W=1u L=180.00n m=1
.ENDS

************************************************************************
* Library Name: VLSI
* Cell Name:    inv
* View Name:    schematic
************************************************************************

.SUBCKT inv IN OUT VDD VSS
*.PININFO IN:I OUT:O VDD:B VSS:B
Mm2 OUT IN VSS VSS n_18 W=500.0n L=180n m=1
Mm1 OUT IN VDD VDD p_18 W=1.85u L=180n m=1
.ENDS

************************************************************************
* Library Name: VLSI
* Cell Name:    DFFTG
* View Name:    schematic
************************************************************************

.SUBCKT DFFTG CLK D Q QM VDD VSS
*.PININFO CLK:I D:B Q:B QM:B VDD:B VSS:B
XI10 net32 net8 CLK net56 VDD VSS / TG
XI9 net36 net8 net56 CLK VDD VSS / TG
XI3 net48 net26 CLK net56 VDD VSS / TG
XI2 net52 net26 net56 CLK VDD VSS / TG
XI13 QM net32 VDD VSS / inv
XI12 Q net36 VDD VSS / inv
XI11 net8 Q VDD VSS / inv
XI5 net26 QM VDD VSS / inv
XI4 QM net48 VDD VSS / inv
XI1 D net52 VDD VSS / inv
XI0 CLK net56 VDD VSS / inv
.ENDS
