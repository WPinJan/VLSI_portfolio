* File: Gal_LFSR.pex.spi
* Created: Thu Dec  5 17:36:50 2024
* Program "Calibre xRC"
* Version "v2016.4_15.11"
* 
.include "Gal_LFSR.pex.spi.pex"
.subckt Gal_LFSR  Q[8] RESET CLK VDD VSS Q[7] Q[1] Q[2] Q[4] Q[5] Q[3] Q[6]
* 
* Q[6]	Q[6]
* Q[3]	Q[3]
* Q[5]	Q[5]
* Q[4]	Q[4]
* Q[2]	Q[2]
* Q[1]	Q[1]
* Q[7]	Q[7]
* VSS	VSS
* VDD	VDD
* CLK	CLK
* RESET	RESET
* Q[8]	Q[8]
mXI16/MM0 N_XI16/NET47_XI16/MM0_d N_Q[4]_XI16/MM0_g N_VSS_XI16/MM0_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI20/MM0 N_XI20/NET47_XI20/MM0_d N_Q[8]_XI20/MM0_g N_VSS_XI20/MM0_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI13/MM3 N_Q[8]_XI13/MM3_d N_NET093_XI13/MM3_g N_VSS_XI13/MM3_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI17/MM3 N_Q[4]_XI17/MM3_d N_QBAR[4]_XI17/MM3_g N_VSS_XI17/MM3_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI16/MM9 N_XI16/NET31_XI16/MM9_d N_XI16/NET47_XI16/MM9_g
+ N_XI16/NET43_XI16/MM9_s N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.125e-13 PD=1.48e-06 PS=8.5e-07
mXI20/MM9 N_XI20/NET31_XI20/MM9_d N_XI20/NET47_XI20/MM9_g
+ N_XI20/NET43_XI20/MM9_s N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.125e-13 PD=1.48e-06 PS=8.5e-07
mXI16/MM1 N_XI16/NET43_XI16/MM1_d N_CLK_XI16/MM1_g N_VSS_XI16/MM1_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.125e-13 AS=2.45e-13 PD=8.5e-07
+ PS=1.48e-06
mXI20/MM1 N_XI20/NET43_XI20/MM1_d N_CLK_XI20/MM1_g N_VSS_XI20/MM1_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.125e-13 AS=2.45e-13 PD=8.5e-07
+ PS=1.48e-06
mXI13/MM2 N_XI13/NET39_XI13/MM2_d N_XI13/NET31_XI13/MM2_g N_VSS_XI13/MM2_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.25e-13 AS=2.45e-13 PD=5e-07
+ PS=1.48e-06
mXI17/MM2 N_XI17/NET39_XI17/MM2_d N_XI17/NET31_XI17/MM2_g N_VSS_XI17/MM2_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.25e-13 AS=2.45e-13 PD=5e-07
+ PS=1.48e-06
mXI13/MM10 N_NET093_XI13/MM10_d N_CLK_XI13/MM10_g N_XI13/NET39_XI13/MM10_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.25e-13 PD=1.48e-06
+ PS=5e-07
mXI17/MM10 N_QBAR[4]_XI17/MM10_d N_CLK_XI17/MM10_g N_XI17/NET39_XI17/MM10_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.25e-13 PD=1.48e-06
+ PS=5e-07
mXI16/MM10 N_QBAR[5]_XI16/MM10_d N_CLK_XI16/MM10_g N_XI16/NET39_XI16/MM10_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.25e-13 PD=1.48e-06
+ PS=5e-07
mXI20/MM10 N_NET0106_XI20/MM10_d N_CLK_XI20/MM10_g N_XI20/NET39_XI20/MM10_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.25e-13 PD=1.48e-06
+ PS=5e-07
mXI16/MM2 N_XI16/NET39_XI16/MM2_d N_XI16/NET31_XI16/MM2_g N_VSS_XI16/MM2_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.25e-13 AS=2.45e-13 PD=5e-07
+ PS=1.48e-06
mXI20/MM2 N_XI20/NET39_XI20/MM2_d N_XI20/NET31_XI20/MM2_g N_VSS_XI20/MM2_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.25e-13 AS=2.45e-13 PD=5e-07
+ PS=1.48e-06
mXI13/MM1 N_XI13/NET43_XI13/MM1_d N_CLK_XI13/MM1_g N_VSS_XI13/MM1_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.125e-13 AS=2.45e-13 PD=8.5e-07
+ PS=1.48e-06
mXI17/MM1 N_XI17/NET43_XI17/MM1_d N_CLK_XI17/MM1_g N_VSS_XI17/MM1_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.125e-13 AS=2.45e-13 PD=8.5e-07
+ PS=1.48e-06
mXI13/MM9 N_XI13/NET31_XI13/MM9_d N_XI13/NET47_XI13/MM9_g
+ N_XI13/NET43_XI13/MM9_s N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.125e-13 PD=1.48e-06 PS=8.5e-07
mXI17/MM9 N_XI17/NET31_XI17/MM9_d N_XI17/NET47_XI17/MM9_g
+ N_XI17/NET43_XI17/MM9_s N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.125e-13 PD=1.48e-06 PS=8.5e-07
mXI16/MM3 N_Q[5]_XI16/MM3_d N_QBAR[5]_XI16/MM3_g N_VSS_XI16/MM3_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI20/MM3 N_Q[1]_XI20/MM3_d N_NET0106_XI20/MM3_g N_VSS_XI20/MM3_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI13/MM0 N_XI13/NET47_XI13/MM0_d N_NET59_XI13/MM0_g N_VSS_XI13/MM0_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI17/MM0 N_XI17/NET47_XI17/MM0_d N_Q[3]_XI17/MM0_g N_VSS_XI17/MM0_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI15/MM0 N_XI15/NET47_XI15/MM0_d N_Q[5]_XI15/MM0_g N_VSS_XI15/MM0_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI8/XI2/MM0 N_NET0113_XI8/XI2/MM0_d N_Q[8]_XI8/XI2/MM0_g N_NET59_XI8/XI2/MM0_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI9/XI3/MM0 N_Q[1]_XI9/XI3/MM0_d N_NET093_XI9/XI3/MM0_g N_NET35_XI9/XI3/MM0_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI18/MM3 N_Q[3]_XI18/MM3_d N_QBAR[3]_XI18/MM3_g N_VSS_XI18/MM3_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI15/MM9 N_XI15/NET31_XI15/MM9_d N_XI15/NET47_XI15/MM9_g
+ N_XI15/NET43_XI15/MM9_s N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.125e-13 PD=1.48e-06 PS=8.5e-07
mXI8/XI3/MM0 N_Q[7]_XI8/XI3/MM0_d N_NET093_XI8/XI3/MM0_g N_NET59_XI8/XI3/MM0_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI9/XI2/MM0 N_NET0106_XI9/XI2/MM0_d N_Q[8]_XI9/XI2/MM0_g N_NET35_XI9/XI2/MM0_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI15/MM1 N_XI15/NET43_XI15/MM1_d N_CLK_XI15/MM1_g N_VSS_XI15/MM1_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.125e-13 AS=2.45e-13 PD=8.5e-07
+ PS=1.48e-06
mXI18/MM2 N_XI18/NET39_XI18/MM2_d N_XI18/NET31_XI18/MM2_g N_VSS_XI18/MM2_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.25e-13 AS=2.45e-13 PD=5e-07
+ PS=1.48e-06
mXI18/MM10 N_QBAR[3]_XI18/MM10_d N_CLK_XI18/MM10_g N_XI18/NET39_XI18/MM10_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.25e-13 PD=1.48e-06
+ PS=5e-07
mXI15/MM10 N_QBAR[6]_XI15/MM10_d N_CLK_XI15/MM10_g N_XI15/NET39_XI15/MM10_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.25e-13 PD=1.48e-06
+ PS=5e-07
mXI19/MM0 N_XI19/NET47_XI19/MM0_d N_NET35_XI19/MM0_g N_VSS_XI19/MM0_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI15/MM2 N_XI15/NET39_XI15/MM2_d N_XI15/NET31_XI15/MM2_g N_VSS_XI15/MM2_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.25e-13 AS=2.45e-13 PD=5e-07
+ PS=1.48e-06
mXI18/MM1 N_XI18/NET43_XI18/MM1_d N_CLK_XI18/MM1_g N_VSS_XI18/MM1_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.125e-13 AS=2.45e-13 PD=8.5e-07
+ PS=1.48e-06
mXI14/MM3 N_Q[7]_XI14/MM3_d N_NET0113_XI14/MM3_g N_VSS_XI14/MM3_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI19/MM9 N_XI19/NET31_XI19/MM9_d N_XI19/NET47_XI19/MM9_g
+ N_XI19/NET43_XI19/MM9_s N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.125e-13 PD=1.48e-06 PS=8.5e-07
mXI18/MM9 N_XI18/NET31_XI18/MM9_d N_XI18/NET47_XI18/MM9_g
+ N_XI18/NET43_XI18/MM9_s N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.125e-13 PD=1.48e-06 PS=8.5e-07
mXI15/MM3 N_Q[6]_XI15/MM3_d N_QBAR[6]_XI15/MM3_g N_VSS_XI15/MM3_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI19/MM1 N_XI19/NET43_XI19/MM1_d N_CLK_XI19/MM1_g N_VSS_XI19/MM1_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.125e-13 AS=2.45e-13 PD=8.5e-07
+ PS=1.48e-06
mXI14/MM2 N_XI14/NET39_XI14/MM2_d N_XI14/NET31_XI14/MM2_g N_VSS_XI14/MM2_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.25e-13 AS=2.45e-13 PD=5e-07
+ PS=1.48e-06
mXI18/MM0 N_XI18/NET47_XI18/MM0_d N_NET23_XI18/MM0_g N_VSS_XI18/MM0_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI14/MM10 N_NET0113_XI14/MM10_d N_CLK_XI14/MM10_g N_XI14/NET39_XI14/MM10_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.25e-13 PD=1.48e-06
+ PS=5e-07
mXI19/MM10 N_NET099_XI19/MM10_d N_CLK_XI19/MM10_g N_XI19/NET39_XI19/MM10_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=1.25e-13 PD=1.48e-06
+ PS=5e-07
mXI19/MM2 N_XI19/NET39_XI19/MM2_d N_XI19/NET31_XI19/MM2_g N_VSS_XI19/MM2_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=1.25e-13 AS=2.45e-13 PD=5e-07
+ PS=1.48e-06
mXI10/XI3/MM0 N_Q[2]_XI10/XI3/MM0_d N_NET093_XI10/XI3/MM0_g
+ N_NET23_XI10/XI3/MM0_s N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI14/MM1 N_XI14/NET43_XI14/MM1_d N_CLK_XI14/MM1_g N_VSS_XI14/MM1_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.125e-13 AS=2.45e-13 PD=8.5e-07
+ PS=1.48e-06
mXI14/MM9 N_XI14/NET31_XI14/MM9_d N_XI14/NET47_XI14/MM9_g
+ N_XI14/NET43_XI14/MM9_s N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.125e-13 PD=1.48e-06 PS=8.5e-07
mXI19/MM3 N_Q[2]_XI19/MM3_d N_NET099_XI19/MM3_g N_VSS_XI19/MM3_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI10/XI2/MM0 N_NET099_XI10/XI2/MM0_d N_Q[8]_XI10/XI2/MM0_g
+ N_NET23_XI10/XI2/MM0_s N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI14/MM0 N_XI14/NET47_XI14/MM0_d N_Q[6]_XI14/MM0_g N_VSS_XI14/MM0_s
+ N_VSS_XI16/MM0_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI13/MM11 N_Q[8]_XI13/MM11_d N_RESET_XI13/MM11_g N_VDD_XI13/MM11_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI16/MM5 N_XI16/NET26_XI16/MM5_d N_Q[4]_XI16/MM5_g N_VDD_XI16/MM5_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=4.59e-13 AS=8.82e-13 PD=5.1e-07
+ PS=2.78e-06
mXI17/MM11 N_Q[4]_XI17/MM11_d N_RESET_XI17/MM11_g N_VDD_XI17/MM11_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI20/MM5 N_XI20/NET26_XI20/MM5_d N_Q[8]_XI20/MM5_g N_VDD_XI20/MM5_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=4.59e-13 AS=8.82e-13 PD=5.1e-07
+ PS=2.78e-06
mXI16/MM4 N_XI16/NET47_XI16/MM4_d N_CLK_XI16/MM4_g N_XI16/NET26_XI16/MM4_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=4.59e-13 PD=2.78e-06
+ PS=5.1e-07
mXI20/MM4 N_XI20/NET47_XI20/MM4_d N_CLK_XI20/MM4_g N_XI20/NET26_XI20/MM4_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=4.59e-13 PD=2.78e-06
+ PS=5.1e-07
mXI13/MM8 N_Q[8]_XI13/MM8_d N_NET093_XI13/MM8_g N_VDD_XI13/MM8_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI17/MM8 N_Q[4]_XI17/MM8_d N_QBAR[4]_XI17/MM8_g N_VDD_XI17/MM8_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI16/MM6 N_XI16/NET31_XI16/MM6_d N_CLK_XI16/MM6_g N_VDD_XI16/MM6_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI20/MM6 N_XI20/NET31_XI20/MM6_d N_CLK_XI20/MM6_g N_VDD_XI20/MM6_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI13/MM7 N_NET093_XI13/MM7_d N_XI13/NET31_XI13/MM7_g N_VDD_XI13/MM7_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI17/MM7 N_QBAR[4]_XI17/MM7_d N_XI17/NET31_XI17/MM7_g N_VDD_XI17/MM7_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI16/MM7 N_QBAR[5]_XI16/MM7_d N_XI16/NET31_XI16/MM7_g N_VDD_XI16/MM7_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI20/MM7 N_NET0106_XI20/MM7_d N_XI20/NET31_XI20/MM7_g N_VDD_XI20/MM7_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI13/MM6 N_XI13/NET31_XI13/MM6_d N_CLK_XI13/MM6_g N_VDD_XI13/MM6_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI17/MM6 N_XI17/NET31_XI17/MM6_d N_CLK_XI17/MM6_g N_VDD_XI17/MM6_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI16/MM8 N_Q[5]_XI16/MM8_d N_QBAR[5]_XI16/MM8_g N_VDD_XI16/MM8_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI20/MM8 N_Q[1]_XI20/MM8_d N_NET0106_XI20/MM8_g N_VDD_XI20/MM8_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI13/MM4 N_XI13/NET47_XI13/MM4_d N_CLK_XI13/MM4_g N_XI13/NET26_XI13/MM4_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=4.59e-13 PD=2.78e-06
+ PS=5.1e-07
mXI17/MM4 N_XI17/NET47_XI17/MM4_d N_CLK_XI17/MM4_g N_XI17/NET26_XI17/MM4_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=4.59e-13 PD=2.78e-06
+ PS=5.1e-07
mXI13/MM5 N_XI13/NET26_XI13/MM5_d N_NET59_XI13/MM5_g N_VDD_XI13/MM5_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=4.59e-13 AS=8.82e-13 PD=5.1e-07
+ PS=2.78e-06
mXI16/MM11 N_Q[5]_XI16/MM11_d N_RESET_XI16/MM11_g N_VDD_XI16/MM11_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI17/MM5 N_XI17/NET26_XI17/MM5_d N_Q[3]_XI17/MM5_g N_VDD_XI17/MM5_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=4.59e-13 AS=8.82e-13 PD=5.1e-07
+ PS=2.78e-06
mXI20/MM11 N_Q[1]_XI20/MM11_d N_RESET_XI20/MM11_g N_VDD_XI20/MM11_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI15/MM5 N_XI15/NET26_XI15/MM5_d N_Q[5]_XI15/MM5_g N_VDD_XI15/MM5_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=4.59e-13 AS=8.82e-13 PD=5.1e-07
+ PS=2.78e-06
mXI18/MM11 N_Q[3]_XI18/MM11_d N_RESET_XI18/MM11_g N_VDD_XI18/MM11_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI8/XI3/MM1 N_Q[7]_XI8/XI3/MM1_d N_Q[8]_XI8/XI3/MM1_g N_NET59_XI8/XI3/MM1_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI9/XI2/MM1 N_NET0106_XI9/XI2/MM1_d N_NET093_XI9/XI2/MM1_g
+ N_NET35_XI9/XI2/MM1_s N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI15/MM4 N_XI15/NET47_XI15/MM4_d N_CLK_XI15/MM4_g N_XI15/NET26_XI15/MM4_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=4.59e-13 PD=2.78e-06
+ PS=5.1e-07
mXI18/MM8 N_Q[3]_XI18/MM8_d N_QBAR[3]_XI18/MM8_g N_VDD_XI18/MM8_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI8/XI2/MM1 N_NET0113_XI8/XI2/MM1_d N_NET093_XI8/XI2/MM1_g
+ N_NET59_XI8/XI2/MM1_s N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI9/XI3/MM1 N_Q[1]_XI9/XI3/MM1_d N_Q[8]_XI9/XI3/MM1_g N_NET35_XI9/XI3/MM1_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI15/MM6 N_XI15/NET31_XI15/MM6_d N_CLK_XI15/MM6_g N_VDD_XI15/MM6_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI18/MM7 N_QBAR[3]_XI18/MM7_d N_XI18/NET31_XI18/MM7_g N_VDD_XI18/MM7_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI14/MM11 N_Q[7]_XI14/MM11_d N_RESET_XI14/MM11_g N_VDD_XI14/MM11_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI19/MM5 N_XI19/NET26_XI19/MM5_d N_NET35_XI19/MM5_g N_VDD_XI19/MM5_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=4.59e-13 AS=8.82e-13 PD=5.1e-07
+ PS=2.78e-06
mXI15/MM7 N_QBAR[6]_XI15/MM7_d N_XI15/NET31_XI15/MM7_g N_VDD_XI15/MM7_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI19/MM4 N_XI19/NET47_XI19/MM4_d N_CLK_XI19/MM4_g N_XI19/NET26_XI19/MM4_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=4.59e-13 PD=2.78e-06
+ PS=5.1e-07
mXI18/MM6 N_XI18/NET31_XI18/MM6_d N_CLK_XI18/MM6_g N_VDD_XI18/MM6_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI14/MM8 N_Q[7]_XI14/MM8_d N_NET0113_XI14/MM8_g N_VDD_XI14/MM8_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI15/MM8 N_Q[6]_XI15/MM8_d N_QBAR[6]_XI15/MM8_g N_VDD_XI15/MM8_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI19/MM6 N_XI19/NET31_XI19/MM6_d N_CLK_XI19/MM6_g N_VDD_XI19/MM6_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI18/MM4 N_XI18/NET47_XI18/MM4_d N_CLK_XI18/MM4_g N_XI18/NET26_XI18/MM4_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=4.59e-13 PD=2.78e-06
+ PS=5.1e-07
mXI14/MM7 N_NET0113_XI14/MM7_d N_XI14/NET31_XI14/MM7_g N_VDD_XI14/MM7_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI15/MM11 N_Q[6]_XI15/MM11_d N_RESET_XI15/MM11_g N_VDD_XI15/MM11_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI18/MM5 N_XI18/NET26_XI18/MM5_d N_NET23_XI18/MM5_g N_VDD_XI18/MM5_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=4.59e-13 AS=8.82e-13 PD=5.1e-07
+ PS=2.78e-06
mXI19/MM7 N_NET099_XI19/MM7_d N_XI19/NET31_XI19/MM7_g N_VDD_XI19/MM7_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI10/XI2/MM1 N_NET099_XI10/XI2/MM1_d N_NET093_XI10/XI2/MM1_g
+ N_NET23_XI10/XI2/MM1_s N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI14/MM6 N_XI14/NET31_XI14/MM6_d N_CLK_XI14/MM6_g N_VDD_XI14/MM6_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI19/MM8 N_Q[2]_XI19/MM8_d N_NET099_XI19/MM8_g N_VDD_XI19/MM8_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
mXI10/XI3/MM1 N_Q[2]_XI10/XI3/MM1_d N_Q[8]_XI10/XI3/MM1_g N_NET23_XI10/XI3/MM1_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13
+ PD=1.45e-06 PS=1.45e-06
mXI14/MM4 N_XI14/NET47_XI14/MM4_d N_CLK_XI14/MM4_g N_XI14/NET26_XI14/MM4_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=4.59e-13 PD=2.78e-06
+ PS=5.1e-07
mXI14/MM5 N_XI14/NET26_XI14/MM5_d N_Q[6]_XI14/MM5_g N_VDD_XI14/MM5_s
+ N_VDD_XI13/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=4.59e-13 AS=8.82e-13 PD=5.1e-07
+ PS=2.78e-06
mXI19/MM11 N_Q[2]_XI19/MM11_d N_RESET_XI19/MM11_g N_VDD_XI19/MM11_s
+ N_VDD_XI17/MM11_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13 AS=8.82e-13 PD=2.78e-06
+ PS=2.78e-06
*
.include "Gal_LFSR.pex.spi.GAL_LFSR.pxi"
*
.ends
*
*
