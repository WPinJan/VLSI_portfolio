* File: DFFnand.pex.spi
* Created: Fri Nov 15 20:54:07 2024
* Program "Calibre xRC"
* Version "v2016.4_15.11"
* 
.include "DFFnand.pex.spi.pex"
.subckt DFFnand  VDD VSS QBAR QM Q D CLK
* 
* CLK	CLK
* D	D
* Q	Q
* QM	QM
* QBAR	QBAR
* VSS	VSS
* VDD	VDD
mXI0/MM0 N_XI0/NET14_XI0/MM0_d N_D_XI0/MM0_g N_VSS_XI0/MM0_s N_VSS_XI0/MM0_b
+ N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI9/Mm2 N_NET9_XI9/Mm2_d N_CLK_XI9/Mm2_g N_VSS_XI9/Mm2_s N_VSS_XI0/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI0/MM1 N_NET47_XI0/MM1_d N_NET9_XI0/MM1_g N_XI0/NET14_XI0/MM1_s
+ N_VSS_XI0/MM0_b N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
mXI2/MM1 N_QM_XI2/MM1_d N_NET41_XI2/MM1_g N_XI2/NET14_XI2/MM1_s N_VSS_XI0/MM0_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
mXI2/MM0 N_XI2/NET14_XI2/MM0_d N_NET47_XI2/MM0_g N_VSS_XI2/MM0_s N_VSS_XI0/MM0_b
+ N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI1/MM1 N_XI1/NET14_XI1/MM1_d N_NET9_XI1/MM1_g N_VSS_XI1/MM1_s N_VSS_XI0/MM0_b
+ N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI3/MM1 N_NET41_XI3/MM1_d N_NET48_XI3/MM1_g N_XI3/NET14_XI3/MM1_s
+ N_VSS_XI0/MM0_b N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
mXI1/MM0 N_NET48_XI1/MM0_d N_NET47_XI1/MM0_g N_XI1/NET14_XI1/MM0_s
+ N_VSS_XI0/MM0_b N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
mXI3/MM0 N_XI3/NET14_XI3/MM0_d N_QM_XI3/MM0_g N_VSS_XI3/MM0_s N_VSS_XI0/MM0_b
+ N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI5/MM1 N_Q_XI5/MM1_d N_QBAR_XI5/MM1_g N_XI5/NET14_XI5/MM1_s N_VSS_XI0/MM0_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06 PS=5.1e-07
mXI5/MM0 N_XI5/NET14_XI5/MM0_d N_NET22_XI5/MM0_g N_VSS_XI5/MM0_s N_VSS_XI0/MM0_b
+ N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI7/MM0 N_XI7/NET14_XI7/MM0_d N_QM_XI7/MM0_g N_VSS_XI7/MM0_s N_VSS_XI0/MM0_b
+ N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI8/Mm2 N_NET13_XI8/Mm2_d N_NET9_XI8/Mm2_g N_VSS_XI8/Mm2_s N_VSS_XI0/MM0_b N_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI7/MM1 N_NET22_XI7/MM1_d N_NET13_XI7/MM1_g N_XI7/NET14_XI7/MM1_s
+ N_VSS_XI0/MM0_b N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
mXI6/MM1 N_XI6/NET14_XI6/MM1_d N_NET13_XI6/MM1_g N_VSS_XI6/MM1_s N_VSS_XI0/MM0_b
+ N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI4/MM1 N_QBAR_XI4/MM1_d N_NET23_XI4/MM1_g N_XI4/NET14_XI4/MM1_s
+ N_VSS_XI0/MM0_b N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
mXI6/MM0 N_NET23_XI6/MM0_d N_NET22_XI6/MM0_g N_XI6/NET14_XI6/MM0_s
+ N_VSS_XI0/MM0_b N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=2.55e-13 PD=1.98e-06
+ PS=5.1e-07
mXI4/MM0 N_XI4/NET14_XI4/MM0_d N_Q_XI4/MM0_g N_VSS_XI4/MM0_s N_VSS_XI0/MM0_b
+ N_18 L=1.8e-07 W=1e-06 AD=2.55e-13 AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI0/MM3 N_NET47_XI0/MM3_d N_D_XI0/MM3_g N_VDD_XI0/MM3_s N_VDD_XI0/MM3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI2/MM2 N_QM_XI2/MM2_d N_NET41_XI2/MM2_g N_VDD_XI2/MM2_s N_VDD_XI0/MM3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI2/MM3 N_QM_XI2/MM3_d N_NET47_XI2/MM3_g N_VDD_XI2/MM3_s N_VDD_XI0/MM3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI9/Mm1 N_NET9_XI9/Mm1_d N_CLK_XI9/Mm1_g N_VDD_XI9/Mm1_s N_VDD_XI9/Mm1_b P_18
+ L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXI0/MM2 N_NET47_XI0/MM2_d N_NET9_XI0/MM2_g N_VDD_XI0/MM2_s N_VDD_XI0/MM3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI1/MM2 N_NET48_XI1/MM2_d N_NET9_XI1/MM2_g N_VDD_XI1/MM2_s N_VDD_XI9/Mm1_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI3/MM2 N_NET41_XI3/MM2_d N_NET48_XI3/MM2_g N_VDD_XI3/MM2_s N_VDD_XI0/MM3_b
+ P_18 L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI1/MM3 N_NET48_XI1/MM3_d N_NET47_XI1/MM3_g N_VDD_XI1/MM3_s N_VDD_XI9/Mm1_b
+ P_18 L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI3/MM3 N_NET41_XI3/MM3_d N_QM_XI3/MM3_g N_VDD_XI3/MM3_s N_VDD_XI0/MM3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI7/MM3 N_NET22_XI7/MM3_d N_QM_XI7/MM3_g N_VDD_XI7/MM3_s N_VDD_XI0/MM3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI8/Mm1 N_NET13_XI8/Mm1_d N_NET9_XI8/Mm1_g N_VDD_XI8/Mm1_s N_VDD_XI9/Mm1_b P_18
+ L=1.8e-07 W=1.85e-06 AD=9.065e-13 AS=9.065e-13 PD=2.83e-06 PS=2.83e-06
mXI7/MM2 N_NET22_XI7/MM2_d N_NET13_XI7/MM2_g N_VDD_XI7/MM2_s N_VDD_XI0/MM3_b
+ P_18 L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI5/MM2 N_Q_XI5/MM2_d N_QBAR_XI5/MM2_g N_VDD_XI5/MM2_s N_VDD_XI0/MM3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI5/MM3 N_Q_XI5/MM3_d N_NET22_XI5/MM3_g N_VDD_XI5/MM3_s N_VDD_XI0/MM3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI6/MM2 N_NET23_XI6/MM2_d N_NET13_XI6/MM2_g N_VDD_XI6/MM2_s N_VDD_XI9/Mm1_b
+ P_18 L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI4/MM2 N_QBAR_XI4/MM2_d N_NET23_XI4/MM2_g N_VDD_XI4/MM2_s N_VDD_XI0/MM3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI6/MM3 N_NET23_XI6/MM3_d N_NET22_XI6/MM3_g N_VDD_XI6/MM3_s N_VDD_XI9/Mm1_b
+ P_18 L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
mXI4/MM3 N_QBAR_XI4/MM3_d N_Q_XI4/MM3_g N_VDD_XI4/MM3_s N_VDD_XI0/MM3_b P_18
+ L=1.8e-07 W=1.85e-06 AD=4.7175e-13 AS=9.065e-13 PD=5.1e-07 PS=2.83e-06
*
.include "DFFnand.pex.spi.DFFNAND.pxi"
*
.ends
*
*
