************************************************************************
* auCdl Netlist:
* 
* Library Name:  VLSI
* Top Cell Name: Gal_LFSR
* View Name:     schematic
* Netlisted on:  Dec  2 15:34:51 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: VLSI
* Cell Name:    DFF_dynamic
* View Name:    schematic
************************************************************************

.SUBCKT DFF_dynamic CLK D Q Qbar VDD VSS reset
*.PININFO CLK:I D:I reset:I Q:O Qbar:O VDD:B VSS:B
MM11 Q reset VDD VDD P_18 W=1.8u L=180.00n m=1
MM8 Q Qbar VDD VDD P_18 W=1.8u L=180.00n m=1
MM7 Qbar net31 VDD VDD P_18 W=1.8u L=180.00n m=1
MM6 net31 CLK VDD VDD P_18 W=1.8u L=180.00n m=1
MM5 net26 D VDD VDD P_18 W=1.8u L=180.00n m=1
MM4 net47 CLK net26 VDD P_18 W=1.8u L=180.00n m=1
MM10 Qbar CLK net39 VSS N_18 W=500.0n L=180.00n m=1
MM9 net31 net47 net43 VSS N_18 W=500.0n L=180.00n m=1
MM3 Q Qbar VSS VSS N_18 W=500.0n L=180.00n m=1
MM2 net39 net31 VSS VSS N_18 W=500.0n L=180.00n m=1
MM1 net43 CLK VSS VSS N_18 W=500.0n L=180.00n m=1
MM0 net47 D VSS VSS N_18 W=500.0n L=180.00n m=1
.ENDS

************************************************************************
* Library Name: VLSI
* Cell Name:    TG
* View Name:    schematic
************************************************************************

.SUBCKT TG A B EN ENbar VDD VSS
*.PININFO EN:I ENbar:I A:B B:B VDD:B VSS:B
MM1 A ENbar B VDD P_18 W=470.00n L=180.00n m=1
MM0 A EN B VSS N_18 W=470.00n L=180.00n m=1
.ENDS

************************************************************************
* Library Name: VLSI
* Cell Name:    XOR
* View Name:    schematic
************************************************************************

.SUBCKT XOR A Abar B Bbar VDD VSS Y
*.PININFO A:I Abar:I B:I Bbar:I Y:O VDD:B VSS:B
XI3 B Y Abar A VDD VSS / TG
XI2 Bbar Y A Abar VDD VSS / TG
.ENDS

************************************************************************
* Library Name: VLSI
* Cell Name:    Gal_LFSR
* View Name:    schematic
************************************************************************

.SUBCKT Gal_LFSR CLK Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] Q[8] VDD VSS reset
*.PININFO CLK:I reset:I Qbar[3]:O Qbar[4]:O Qbar[5]:O Qbar[6]:O Q[1]:B Q[2]:B 
*.PININFO Q[3]:B Q[4]:B Q[5]:B Q[6]:B Q[7]:B Q[8]:B VDD:B VSS:B
XI15 CLK Q[5] Q[6] Qbar[6] VDD VSS reset / DFF_dynamic
XI14 CLK Q[6] Q[7] net0113 VDD VSS reset / DFF_dynamic
XI20 CLK Q[8] Q[1] net0106 VDD VSS reset / DFF_dynamic
XI18 CLK net23 Q[3] Qbar[3] VDD VSS reset / DFF_dynamic
XI17 CLK Q[3] Q[4] Qbar[4] VDD VSS reset / DFF_dynamic
XI16 CLK Q[4] Q[5] Qbar[5] VDD VSS reset / DFF_dynamic
XI19 CLK net35 Q[2] net099 VDD VSS reset / DFF_dynamic
XI13 CLK net59 Q[8] net093 VDD VSS reset / DFF_dynamic
XI10 Q[8] net093 Q[2] net099 VDD VSS net23 / XOR
XI9 Q[8] net093 Q[1] net0106 VDD VSS net35 / XOR
XI8 Q[8] net093 Q[7] net0113 VDD VSS net59 / XOR
.ENDS

