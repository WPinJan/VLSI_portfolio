* File: TBC.pex.spi
* Created: Wed Nov  6 16:01:42 2024
* Program "Calibre xRC"
* Version "v2016.4_15.11"
* 
.include "TBC.pex.spi.pex"
.subckt TBC  VDD VSS T[0] T[1] T[2] T[3] T[4] T[5] T[6] T[7] T[8] T[9] T[10] T[11] T[12]
+ T[13] T[14] B[0] B[1] B[2] B[3]
* 
* T[14]	T[14]
* T[13]	T[13]
* T[12]	T[12]
* T[11]	T[11]
* T[10]	T[10]
* T[9]	T[9]
* T[8]	T[8]
* T[4]	T[4]
* T[5]	T[5]
* T[7]	T[7]
* T[6]	T[6]
* T[3]	T[3]
* T[2]	T[2]
* T[1]	T[1]
* T[0]	T[0]
* B[3]	B[3]
* B[2]	B[2]
* B[1]	B[1]
* B[0]	B[0]
* VDD	VDD
* VSS	VSS
mXI01/MM1 N_XI01/NET14_XI01/MM1_d N_T[0]_XI01/MM1_g N_VSS_XI01/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=8.466e-13 AS=1.6268e-12
+ PD=5.1e-07 PS=4.3e-06
mXInd4/MM3 N_XIND4/NET24_XInd4/MM3_d N_ND13_XInd4/MM3_g N_VSS_XInd4/MM3_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.548e-05 AD=3.9474e-12 AS=7.5852e-12
+ PD=5.1e-07 PS=1.646e-05
mXI01/MM0 N_ND01_XI01/MM0_d N_INV1_XI01/MM0_g N_XI01/NET14_XI01/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=1.6268e-12 AS=8.466e-13
+ PD=4.3e-06 PS=5.1e-07
mXInd4/MM2 N_XIND4/NET28_XInd4/MM2_d N_ND57_XInd4/MM2_g
+ N_XIND4/NET24_XInd4/MM2_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.548e-05
+ AD=3.9474e-12 AS=3.9474e-12 PD=5.1e-07 PS=5.1e-07
mXInd4/MM1 N_XIND4/NET32_XInd4/MM1_d N_ND911_XInd4/MM1_g
+ N_XIND4/NET28_XInd4/MM1_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.548e-05
+ AD=3.9474e-12 AS=3.9474e-12 PD=5.1e-07 PS=5.1e-07
mXInd4/MM0 N_NETB1_XInd4/MM0_d N_INV13_XInd4/MM0_g N_XIND4/NET32_XInd4/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.548e-05 AD=7.5852e-12 AS=3.9474e-12
+ PD=1.646e-05 PS=5.1e-07
mXI1/Mm2 N_INV1_XI1/Mm2_d N_T[1]_XI1/Mm2_g N_VSS_XI1/Mm2_s N_VSS_XI01/MM1_b N_18
+ L=1.8e-07 W=2.08e-06 AD=1.0192e-12 AS=1.0192e-12 PD=3.06e-06 PS=3.06e-06
mXInd22/MM0 N_XIND22/NET14_XInd22/MM0_d N_ND37_XInd22/MM0_g N_VSS_XInd22/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.084e-05 AD=2.7642e-12 AS=5.3116e-12
+ PD=5.1e-07 PS=1.182e-05
mXInd22/MM1 N_NETB2_XInd22/MM1_d N_INV11_XInd22/MM1_g
+ N_XIND22/NET14_XInd22/MM1_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.084e-05
+ AD=5.3116e-12 AS=2.7642e-12 PD=1.182e-05 PS=5.1e-07
mXInd13/MM1 N_XIND13/NET14_XInd13/MM1_d N_T[1]_XInd13/MM1_g N_VSS_XInd13/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=8.466e-13 AS=1.6268e-12
+ PD=5.1e-07 PS=4.3e-06
mXInd13/MM0 N_ND13_XInd13/MM0_d N_INV3_XInd13/MM0_g N_XIND13/NET14_XInd13/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=1.6268e-12 AS=8.466e-13
+ PD=4.3e-06 PS=5.1e-07
mXInd8/MM7 N_XIND8/NET44_XInd8/MM7_d N_INV14_XInd8/MM7_g N_VSS_XInd8/MM7_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.97e-05 AD=5.0235e-12 AS=9.653e-12
+ PD=5.1e-07 PS=2.068e-05
mXInd8/MM6 N_XIND8/NET48_XInd8/MM6_d N_ND67_XInd8/MM6_g
+ N_XIND8/NET44_XInd8/MM6_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.97e-05
+ AD=5.0235e-12 AS=5.0235e-12 PD=5.1e-07 PS=5.1e-07
mXI23/MM1 N_XI23/NET14_XI23/MM1_d N_T[2]_XI23/MM1_g N_VSS_XI23/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=8.466e-13 AS=1.6268e-12
+ PD=5.1e-07 PS=4.3e-06
mXInd8/MM5 N_XIND8/NET52_XInd8/MM5_d N_ND01_XInd8/MM5_g
+ N_XIND8/NET48_XInd8/MM5_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.97e-05
+ AD=5.0235e-12 AS=5.0235e-12 PD=5.1e-07 PS=5.1e-07
mXI23/MM0 N_ND23_XI23/MM0_d N_INV3_XI23/MM0_g N_XI23/NET14_XI23/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=1.6268e-12 AS=8.466e-13
+ PD=4.3e-06 PS=5.1e-07
mXInd8/MM4 N_XIND8/NET56_XInd8/MM4_d N_ND23_XInd8/MM4_g
+ N_XIND8/NET52_XInd8/MM4_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.97e-05
+ AD=5.0235e-12 AS=5.0235e-12 PD=5.1e-07 PS=5.1e-07
mXInd8/MM3 N_XIND8/NET60_XInd8/MM3_d N_ND45_XInd8/MM3_g
+ N_XIND8/NET56_XInd8/MM3_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.97e-05
+ AD=5.0235e-12 AS=5.0235e-12 PD=5.1e-07 PS=5.1e-07
mXInd8/MM2 N_XIND8/NET64_XInd8/MM2_d N_ND89_XInd8/MM2_g
+ N_XIND8/NET60_XInd8/MM2_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.97e-05
+ AD=5.0235e-12 AS=5.0235e-12 PD=5.1e-07 PS=5.1e-07
mXI3/Mm2 N_INV3_XI3/Mm2_d N_T[3]_XI3/Mm2_g N_VSS_XI3/Mm2_s N_VSS_XI01/MM1_b N_18
+ L=1.8e-07 W=2.08e-06 AD=1.0192e-12 AS=1.0192e-12 PD=3.06e-06 PS=3.06e-06
mXInd8/MM0 N_XIND8/NET68_XInd8/MM0_d N_ND1011_XInd8/MM0_g
+ N_XIND8/NET64_XInd8/MM0_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.97e-05
+ AD=5.0235e-12 AS=5.0235e-12 PD=5.1e-07 PS=5.1e-07
mXInd8/MM1 N_NETB0_XInd8/MM1_d N_ND1213_XInd8/MM1_g N_XIND8/NET68_XInd8/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.97e-05 AD=9.653e-12 AS=5.0235e-12
+ PD=2.068e-05 PS=5.1e-07
mXI37/MM1 N_XI37/NET14_XI37/MM1_d N_T[3]_XI37/MM1_g N_VSS_XI37/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=8.466e-13 AS=1.6268e-12
+ PD=5.1e-07 PS=4.3e-06
mXI37/MM0 N_ND37_XI37/MM0_d N_INV7_XI37/MM0_g N_XI37/NET14_XI37/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=1.6268e-12 AS=8.466e-13
+ PD=4.3e-06 PS=5.1e-07
mXIbf0/MM1 N_B[0]_XIbf0/MM1_d N_XIBF0/NET17_XIbf0/MM1_g N_VSS_XIbf0/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07
+ PS=2.48e-06
mXIbf0/MM1@28 N_B[0]_XIbf0/MM1@28_d N_XIBF0/NET17_XIbf0/MM1@28_g
+ N_VSS_XIbf0/MM1@28_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@27 N_B[0]_XIbf0/MM1@27_d N_XIBF0/NET17_XIbf0/MM1@27_g
+ N_VSS_XIbf0/MM1@27_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@26 N_B[0]_XIbf0/MM1@26_d N_XIBF0/NET17_XIbf0/MM1@26_g
+ N_VSS_XIbf0/MM1@26_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@25 N_B[0]_XIbf0/MM1@25_d N_XIBF0/NET17_XIbf0/MM1@25_g
+ N_VSS_XIbf0/MM1@25_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@24 N_B[0]_XIbf0/MM1@24_d N_XIBF0/NET17_XIbf0/MM1@24_g
+ N_VSS_XIbf0/MM1@24_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@23 N_B[0]_XIbf0/MM1@23_d N_XIBF0/NET17_XIbf0/MM1@23_g
+ N_VSS_XIbf0/MM1@23_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@22 N_B[0]_XIbf0/MM1@22_d N_XIBF0/NET17_XIbf0/MM1@22_g
+ N_VSS_XIbf0/MM1@22_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@21 N_B[0]_XIbf0/MM1@21_d N_XIBF0/NET17_XIbf0/MM1@21_g
+ N_VSS_XIbf0/MM1@21_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@20 N_B[0]_XIbf0/MM1@20_d N_XIBF0/NET17_XIbf0/MM1@20_g
+ N_VSS_XIbf0/MM1@20_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@19 N_B[0]_XIbf0/MM1@19_d N_XIBF0/NET17_XIbf0/MM1@19_g
+ N_VSS_XIbf0/MM1@19_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@18 N_B[0]_XIbf0/MM1@18_d N_XIBF0/NET17_XIbf0/MM1@18_g
+ N_VSS_XIbf0/MM1@18_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@17 N_B[0]_XIbf0/MM1@17_d N_XIBF0/NET17_XIbf0/MM1@17_g
+ N_VSS_XIbf0/MM1@17_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@16 N_B[0]_XIbf0/MM1@16_d N_XIBF0/NET17_XIbf0/MM1@16_g
+ N_VSS_XIbf0/MM1@16_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@15 N_B[0]_XIbf0/MM1@15_d N_XIBF0/NET17_XIbf0/MM1@15_g
+ N_VSS_XIbf0/MM1@15_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@14 N_B[0]_XIbf0/MM1@14_d N_XIBF0/NET17_XIbf0/MM1@14_g
+ N_VSS_XIbf0/MM1@14_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@13 N_B[0]_XIbf0/MM1@13_d N_XIBF0/NET17_XIbf0/MM1@13_g
+ N_VSS_XIbf0/MM1@13_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@12 N_B[0]_XIbf0/MM1@12_d N_XIBF0/NET17_XIbf0/MM1@12_g
+ N_VSS_XIbf0/MM1@12_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@11 N_B[0]_XIbf0/MM1@11_d N_XIBF0/NET17_XIbf0/MM1@11_g
+ N_VSS_XIbf0/MM1@11_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@10 N_B[0]_XIbf0/MM1@10_d N_XIBF0/NET17_XIbf0/MM1@10_g
+ N_VSS_XIbf0/MM1@10_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@9 N_B[0]_XIbf0/MM1@9_d N_XIBF0/NET17_XIbf0/MM1@9_g
+ N_VSS_XIbf0/MM1@9_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@8 N_B[0]_XIbf0/MM1@8_d N_XIBF0/NET17_XIbf0/MM1@8_g
+ N_VSS_XIbf0/MM1@8_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@7 N_B[0]_XIbf0/MM1@7_d N_XIBF0/NET17_XIbf0/MM1@7_g
+ N_VSS_XIbf0/MM1@7_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@6 N_B[0]_XIbf0/MM1@6_d N_XIBF0/NET17_XIbf0/MM1@6_g
+ N_VSS_XIbf0/MM1@6_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@5 N_B[0]_XIbf0/MM1@5_d N_XIBF0/NET17_XIbf0/MM1@5_g
+ N_VSS_XIbf0/MM1@5_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@4 N_B[0]_XIbf0/MM1@4_d N_XIBF0/NET17_XIbf0/MM1@4_g
+ N_VSS_XIbf0/MM1@4_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@3 N_B[0]_XIbf0/MM1@3_d N_XIBF0/NET17_XIbf0/MM1@3_g
+ N_VSS_XIbf0/MM1@3_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM1@2 N_B[0]_XIbf0/MM1@2_d N_XIBF0/NET17_XIbf0/MM1@2_g
+ N_VSS_XIbf0/MM1@2_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mXIbf0/MM0 N_XIBF0/NET17_XIbf0/MM0_d N_NETB0_XIbf0/MM0_g N_VSS_XIbf0/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06
+ PS=5.1e-07
mXIbf0/MM0@7 N_XIBF0/NET17_XIbf0/MM0@7_d N_NETB0_XIbf0/MM0@7_g
+ N_VSS_XIbf0/MM0@7_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM0@6 N_XIBF0/NET17_XIbf0/MM0@6_d N_NETB0_XIbf0/MM0@6_g
+ N_VSS_XIbf0/MM0@6_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM0@5 N_XIBF0/NET17_XIbf0/MM0@5_d N_NETB0_XIbf0/MM0@5_g
+ N_VSS_XIbf0/MM0@5_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM0@4 N_XIBF0/NET17_XIbf0/MM0@4_d N_NETB0_XIbf0/MM0@4_g
+ N_VSS_XIbf0/MM0@4_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM0@3 N_XIBF0/NET17_XIbf0/MM0@3_d N_NETB0_XIbf0/MM0@3_g
+ N_VSS_XIbf0/MM0@3_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM0@2 N_XIBF0/NET17_XIbf0/MM0@2_d N_NETB0_XIbf0/MM0@2_g
+ N_VSS_XIbf0/MM0@2_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mXI67/MM1 N_XI67/NET14_XI67/MM1_d N_T[6]_XI67/MM1_g N_VSS_XI67/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=8.466e-13 AS=1.6268e-12
+ PD=5.1e-07 PS=4.3e-06
mXI67/MM0 N_ND67_XI67/MM0_d N_INV7_XI67/MM0_g N_XI67/NET14_XI67/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=1.6268e-12 AS=8.466e-13
+ PD=4.3e-06 PS=5.1e-07
mXIb31/Mm2 N_NETB31_XIb31/Mm2_d N_INV7_XIb31/Mm2_g N_VSS_XIb31/Mm2_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=2.08e-06 AD=1.0192e-12 AS=1.0192e-12
+ PD=3.06e-06 PS=3.06e-06
mXI7/Mm2 N_INV7_XI7/Mm2_d N_T[7]_XI7/Mm2_g N_VSS_XI7/Mm2_s N_VSS_XI01/MM1_b N_18
+ L=1.8e-07 W=2.08e-06 AD=1.0192e-12 AS=1.0192e-12 PD=3.06e-06 PS=3.06e-06
mXI57/MM0 N_XI57/NET14_XI57/MM0_d N_INV7_XI57/MM0_g N_VSS_XI57/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=8.466e-13 AS=1.6268e-12
+ PD=5.1e-07 PS=4.3e-06
mXI57/MM1 N_ND57_XI57/MM1_d N_T[5]_XI57/MM1_g N_XI57/NET14_XI57/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=1.6268e-12 AS=8.466e-13
+ PD=4.3e-06 PS=5.1e-07
mXI5/Mm2 N_INV5_XI5/Mm2_d N_T[5]_XI5/Mm2_g N_VSS_XI5/Mm2_s N_VSS_XI01/MM1_b N_18
+ L=1.8e-07 W=2.08e-06 AD=1.0192e-12 AS=1.0192e-12 PD=3.06e-06 PS=3.06e-06
mXI45/MM0 N_ND45_XI45/MM0_d N_INV5_XI45/MM0_g N_XI45/NET14_XI45/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=1.6268e-12 AS=8.466e-13
+ PD=4.3e-06 PS=5.1e-07
mXI45/MM1 N_XI45/NET14_XI45/MM1_d N_T[4]_XI45/MM1_g N_VSS_XI45/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=8.466e-13 AS=1.6268e-12
+ PD=5.1e-07 PS=4.3e-06
mXIbf1/MM1 N_B[1]_XIbf1/MM1_d N_XIBF1/NET17_XIbf1/MM1_g N_VSS_XIbf1/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07
+ PS=2.48e-06
mXIbf1/MM1@28 N_B[1]_XIbf1/MM1@28_d N_XIBF1/NET17_XIbf1/MM1@28_g
+ N_VSS_XIbf1/MM1@28_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@27 N_B[1]_XIbf1/MM1@27_d N_XIBF1/NET17_XIbf1/MM1@27_g
+ N_VSS_XIbf1/MM1@27_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@26 N_B[1]_XIbf1/MM1@26_d N_XIBF1/NET17_XIbf1/MM1@26_g
+ N_VSS_XIbf1/MM1@26_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@25 N_B[1]_XIbf1/MM1@25_d N_XIBF1/NET17_XIbf1/MM1@25_g
+ N_VSS_XIbf1/MM1@25_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@24 N_B[1]_XIbf1/MM1@24_d N_XIBF1/NET17_XIbf1/MM1@24_g
+ N_VSS_XIbf1/MM1@24_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@23 N_B[1]_XIbf1/MM1@23_d N_XIBF1/NET17_XIbf1/MM1@23_g
+ N_VSS_XIbf1/MM1@23_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@22 N_B[1]_XIbf1/MM1@22_d N_XIBF1/NET17_XIbf1/MM1@22_g
+ N_VSS_XIbf1/MM1@22_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@21 N_B[1]_XIbf1/MM1@21_d N_XIBF1/NET17_XIbf1/MM1@21_g
+ N_VSS_XIbf1/MM1@21_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@20 N_B[1]_XIbf1/MM1@20_d N_XIBF1/NET17_XIbf1/MM1@20_g
+ N_VSS_XIbf1/MM1@20_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@19 N_B[1]_XIbf1/MM1@19_d N_XIBF1/NET17_XIbf1/MM1@19_g
+ N_VSS_XIbf1/MM1@19_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@18 N_B[1]_XIbf1/MM1@18_d N_XIBF1/NET17_XIbf1/MM1@18_g
+ N_VSS_XIbf1/MM1@18_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@17 N_B[1]_XIbf1/MM1@17_d N_XIBF1/NET17_XIbf1/MM1@17_g
+ N_VSS_XIbf1/MM1@17_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@16 N_B[1]_XIbf1/MM1@16_d N_XIBF1/NET17_XIbf1/MM1@16_g
+ N_VSS_XIbf1/MM1@16_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@15 N_B[1]_XIbf1/MM1@15_d N_XIBF1/NET17_XIbf1/MM1@15_g
+ N_VSS_XIbf1/MM1@15_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@14 N_B[1]_XIbf1/MM1@14_d N_XIBF1/NET17_XIbf1/MM1@14_g
+ N_VSS_XIbf1/MM1@14_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@13 N_B[1]_XIbf1/MM1@13_d N_XIBF1/NET17_XIbf1/MM1@13_g
+ N_VSS_XIbf1/MM1@13_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@12 N_B[1]_XIbf1/MM1@12_d N_XIBF1/NET17_XIbf1/MM1@12_g
+ N_VSS_XIbf1/MM1@12_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@11 N_B[1]_XIbf1/MM1@11_d N_XIBF1/NET17_XIbf1/MM1@11_g
+ N_VSS_XIbf1/MM1@11_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@10 N_B[1]_XIbf1/MM1@10_d N_XIBF1/NET17_XIbf1/MM1@10_g
+ N_VSS_XIbf1/MM1@10_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@9 N_B[1]_XIbf1/MM1@9_d N_XIBF1/NET17_XIbf1/MM1@9_g
+ N_VSS_XIbf1/MM1@9_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@8 N_B[1]_XIbf1/MM1@8_d N_XIBF1/NET17_XIbf1/MM1@8_g
+ N_VSS_XIbf1/MM1@8_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@7 N_B[1]_XIbf1/MM1@7_d N_XIBF1/NET17_XIbf1/MM1@7_g
+ N_VSS_XIbf1/MM1@7_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@6 N_B[1]_XIbf1/MM1@6_d N_XIBF1/NET17_XIbf1/MM1@6_g
+ N_VSS_XIbf1/MM1@6_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@5 N_B[1]_XIbf1/MM1@5_d N_XIBF1/NET17_XIbf1/MM1@5_g
+ N_VSS_XIbf1/MM1@5_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@4 N_B[1]_XIbf1/MM1@4_d N_XIBF1/NET17_XIbf1/MM1@4_g
+ N_VSS_XIbf1/MM1@4_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@3 N_B[1]_XIbf1/MM1@3_d N_XIBF1/NET17_XIbf1/MM1@3_g
+ N_VSS_XIbf1/MM1@3_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM1@2 N_B[1]_XIbf1/MM1@2_d N_XIBF1/NET17_XIbf1/MM1@2_g
+ N_VSS_XIbf1/MM1@2_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mXIbf1/MM0 N_XIBF1/NET17_XIbf1/MM0_d N_NETB1_XIbf1/MM0_g N_VSS_XIbf1/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06
+ PS=5.1e-07
mXIbf1/MM0@7 N_XIBF1/NET17_XIbf1/MM0@7_d N_NETB1_XIbf1/MM0@7_g
+ N_VSS_XIbf1/MM0@7_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM0@6 N_XIBF1/NET17_XIbf1/MM0@6_d N_NETB1_XIbf1/MM0@6_g
+ N_VSS_XIbf1/MM0@6_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM0@5 N_XIBF1/NET17_XIbf1/MM0@5_d N_NETB1_XIbf1/MM0@5_g
+ N_VSS_XIbf1/MM0@5_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM0@4 N_XIBF1/NET17_XIbf1/MM0@4_d N_NETB1_XIbf1/MM0@4_g
+ N_VSS_XIbf1/MM0@4_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM0@3 N_XIBF1/NET17_XIbf1/MM0@3_d N_NETB1_XIbf1/MM0@3_g
+ N_VSS_XIbf1/MM0@3_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM0@2 N_XIBF1/NET17_XIbf1/MM0@2_d N_NETB1_XIbf1/MM0@2_g
+ N_VSS_XIbf1/MM0@2_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mXI89/MM1 N_XI89/NET14_XI89/MM1_d N_T[8]_XI89/MM1_g N_VSS_XI89/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=8.466e-13 AS=1.6268e-12
+ PD=5.1e-07 PS=4.3e-06
mXI89/MM0 N_ND89_XI89/MM0_d N_INV9_XI89/MM0_g N_XI89/NET14_XI89/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=1.6268e-12 AS=8.466e-13
+ PD=4.3e-06 PS=5.1e-07
mXIbf2/MM1 N_B[2]_XIbf2/MM1_d N_XIBF2/NET17_XIbf2/MM1_g N_VSS_XIbf2/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07
+ PS=2.48e-06
mXIbf2/MM1@28 N_B[2]_XIbf2/MM1@28_d N_XIBF2/NET17_XIbf2/MM1@28_g
+ N_VSS_XIbf2/MM1@28_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@27 N_B[2]_XIbf2/MM1@27_d N_XIBF2/NET17_XIbf2/MM1@27_g
+ N_VSS_XIbf2/MM1@27_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@26 N_B[2]_XIbf2/MM1@26_d N_XIBF2/NET17_XIbf2/MM1@26_g
+ N_VSS_XIbf2/MM1@26_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@25 N_B[2]_XIbf2/MM1@25_d N_XIBF2/NET17_XIbf2/MM1@25_g
+ N_VSS_XIbf2/MM1@25_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@24 N_B[2]_XIbf2/MM1@24_d N_XIBF2/NET17_XIbf2/MM1@24_g
+ N_VSS_XIbf2/MM1@24_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@23 N_B[2]_XIbf2/MM1@23_d N_XIBF2/NET17_XIbf2/MM1@23_g
+ N_VSS_XIbf2/MM1@23_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@22 N_B[2]_XIbf2/MM1@22_d N_XIBF2/NET17_XIbf2/MM1@22_g
+ N_VSS_XIbf2/MM1@22_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@21 N_B[2]_XIbf2/MM1@21_d N_XIBF2/NET17_XIbf2/MM1@21_g
+ N_VSS_XIbf2/MM1@21_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@20 N_B[2]_XIbf2/MM1@20_d N_XIBF2/NET17_XIbf2/MM1@20_g
+ N_VSS_XIbf2/MM1@20_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@19 N_B[2]_XIbf2/MM1@19_d N_XIBF2/NET17_XIbf2/MM1@19_g
+ N_VSS_XIbf2/MM1@19_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@18 N_B[2]_XIbf2/MM1@18_d N_XIBF2/NET17_XIbf2/MM1@18_g
+ N_VSS_XIbf2/MM1@18_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@17 N_B[2]_XIbf2/MM1@17_d N_XIBF2/NET17_XIbf2/MM1@17_g
+ N_VSS_XIbf2/MM1@17_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@16 N_B[2]_XIbf2/MM1@16_d N_XIBF2/NET17_XIbf2/MM1@16_g
+ N_VSS_XIbf2/MM1@16_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@15 N_B[2]_XIbf2/MM1@15_d N_XIBF2/NET17_XIbf2/MM1@15_g
+ N_VSS_XIbf2/MM1@15_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@14 N_B[2]_XIbf2/MM1@14_d N_XIBF2/NET17_XIbf2/MM1@14_g
+ N_VSS_XIbf2/MM1@14_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@13 N_B[2]_XIbf2/MM1@13_d N_XIBF2/NET17_XIbf2/MM1@13_g
+ N_VSS_XIbf2/MM1@13_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@12 N_B[2]_XIbf2/MM1@12_d N_XIBF2/NET17_XIbf2/MM1@12_g
+ N_VSS_XIbf2/MM1@12_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@11 N_B[2]_XIbf2/MM1@11_d N_XIBF2/NET17_XIbf2/MM1@11_g
+ N_VSS_XIbf2/MM1@11_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@10 N_B[2]_XIbf2/MM1@10_d N_XIBF2/NET17_XIbf2/MM1@10_g
+ N_VSS_XIbf2/MM1@10_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@9 N_B[2]_XIbf2/MM1@9_d N_XIBF2/NET17_XIbf2/MM1@9_g
+ N_VSS_XIbf2/MM1@9_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@8 N_B[2]_XIbf2/MM1@8_d N_XIBF2/NET17_XIbf2/MM1@8_g
+ N_VSS_XIbf2/MM1@8_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@7 N_B[2]_XIbf2/MM1@7_d N_XIBF2/NET17_XIbf2/MM1@7_g
+ N_VSS_XIbf2/MM1@7_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@6 N_B[2]_XIbf2/MM1@6_d N_XIBF2/NET17_XIbf2/MM1@6_g
+ N_VSS_XIbf2/MM1@6_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@5 N_B[2]_XIbf2/MM1@5_d N_XIBF2/NET17_XIbf2/MM1@5_g
+ N_VSS_XIbf2/MM1@5_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@4 N_B[2]_XIbf2/MM1@4_d N_XIBF2/NET17_XIbf2/MM1@4_g
+ N_VSS_XIbf2/MM1@4_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@3 N_B[2]_XIbf2/MM1@3_d N_XIBF2/NET17_XIbf2/MM1@3_g
+ N_VSS_XIbf2/MM1@3_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM1@2 N_B[2]_XIbf2/MM1@2_d N_XIBF2/NET17_XIbf2/MM1@2_g
+ N_VSS_XIbf2/MM1@2_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mXIbf2/MM0 N_XIBF2/NET17_XIbf2/MM0_d N_NETB2_XIbf2/MM0_g N_VSS_XIbf2/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06
+ PS=5.1e-07
mXIbf2/MM0@7 N_XIBF2/NET17_XIbf2/MM0@7_d N_NETB2_XIbf2/MM0@7_g
+ N_VSS_XIbf2/MM0@7_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM0@6 N_XIBF2/NET17_XIbf2/MM0@6_d N_NETB2_XIbf2/MM0@6_g
+ N_VSS_XIbf2/MM0@6_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM0@5 N_XIBF2/NET17_XIbf2/MM0@5_d N_NETB2_XIbf2/MM0@5_g
+ N_VSS_XIbf2/MM0@5_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM0@4 N_XIBF2/NET17_XIbf2/MM0@4_d N_NETB2_XIbf2/MM0@4_g
+ N_VSS_XIbf2/MM0@4_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM0@3 N_XIBF2/NET17_XIbf2/MM0@3_d N_NETB2_XIbf2/MM0@3_g
+ N_VSS_XIbf2/MM0@3_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM0@2 N_XIBF2/NET17_XIbf2/MM0@2_d N_NETB2_XIbf2/MM0@2_g
+ N_VSS_XIbf2/MM0@2_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mXI9/Mm2 N_INV9_XI9/Mm2_d N_T[9]_XI9/Mm2_g N_VSS_XI9/Mm2_s N_VSS_XI01/MM1_b N_18
+ L=1.8e-07 W=2.08e-06 AD=1.0192e-12 AS=1.0192e-12 PD=3.06e-06 PS=3.06e-06
mXI911/MM1 N_XI911/NET14_XI911/MM1_d N_T[9]_XI911/MM1_g N_VSS_XI911/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=8.466e-13 AS=1.6268e-12
+ PD=5.1e-07 PS=4.3e-06
mXI911/MM0 N_ND911_XI911/MM0_d N_INV11_XI911/MM0_g N_XI911/NET14_XI911/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=1.6268e-12 AS=8.466e-13
+ PD=4.3e-06 PS=5.1e-07
mXI1011/MM1 N_XI1011/NET14_XI1011/MM1_d N_T[10]_XI1011/MM1_g N_VSS_XI1011/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=8.466e-13 AS=1.6268e-12
+ PD=5.1e-07 PS=4.3e-06
mXI1011/MM0 N_ND1011_XI1011/MM0_d N_INV11_XI1011/MM0_g
+ N_XI1011/NET14_XI1011/MM0_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06
+ AD=1.6268e-12 AS=8.466e-13 PD=4.3e-06 PS=5.1e-07
mXI11/Mm2 N_INV11_XI11/Mm2_d N_T[11]_XI11/Mm2_g N_VSS_XI11/Mm2_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=2.08e-06 AD=1.0192e-12 AS=1.0192e-12
+ PD=3.06e-06 PS=3.06e-06
mXI1213/MM1 N_XI1213/NET14_XI1213/MM1_d N_T[12]_XI1213/MM1_g N_VSS_XI1213/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06 AD=8.466e-13 AS=1.6268e-12
+ PD=5.1e-07 PS=4.3e-06
mXI1213/MM0 N_ND1213_XI1213/MM0_d N_INV13_XI1213/MM0_g
+ N_XI1213/NET14_XI1213/MM0_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=3.32e-06
+ AD=1.6268e-12 AS=8.466e-13 PD=4.3e-06 PS=5.1e-07
mXI13/Mm2 N_INV13_XI13/Mm2_d N_T[13]_XI13/Mm2_g N_VSS_XI13/Mm2_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=2.08e-06 AD=1.0192e-12 AS=1.0192e-12
+ PD=3.06e-06 PS=3.06e-06
mXIbf3/MM1 N_B[3]_XIbf3/MM1_d N_XIBF3/NET17_XIbf3/MM1_g N_VSS_XIbf3/MM1_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13 AS=7.35e-13 PD=5.1e-07
+ PS=2.48e-06
mXIbf3/MM1@28 N_B[3]_XIbf3/MM1@28_d N_XIBF3/NET17_XIbf3/MM1@28_g
+ N_VSS_XIbf3/MM1@28_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@27 N_B[3]_XIbf3/MM1@27_d N_XIBF3/NET17_XIbf3/MM1@27_g
+ N_VSS_XIbf3/MM1@27_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@26 N_B[3]_XIbf3/MM1@26_d N_XIBF3/NET17_XIbf3/MM1@26_g
+ N_VSS_XIbf3/MM1@26_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@25 N_B[3]_XIbf3/MM1@25_d N_XIBF3/NET17_XIbf3/MM1@25_g
+ N_VSS_XIbf3/MM1@25_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@24 N_B[3]_XIbf3/MM1@24_d N_XIBF3/NET17_XIbf3/MM1@24_g
+ N_VSS_XIbf3/MM1@24_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@23 N_B[3]_XIbf3/MM1@23_d N_XIBF3/NET17_XIbf3/MM1@23_g
+ N_VSS_XIbf3/MM1@23_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@22 N_B[3]_XIbf3/MM1@22_d N_XIBF3/NET17_XIbf3/MM1@22_g
+ N_VSS_XIbf3/MM1@22_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@21 N_B[3]_XIbf3/MM1@21_d N_XIBF3/NET17_XIbf3/MM1@21_g
+ N_VSS_XIbf3/MM1@21_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@20 N_B[3]_XIbf3/MM1@20_d N_XIBF3/NET17_XIbf3/MM1@20_g
+ N_VSS_XIbf3/MM1@20_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@19 N_B[3]_XIbf3/MM1@19_d N_XIBF3/NET17_XIbf3/MM1@19_g
+ N_VSS_XIbf3/MM1@19_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@18 N_B[3]_XIbf3/MM1@18_d N_XIBF3/NET17_XIbf3/MM1@18_g
+ N_VSS_XIbf3/MM1@18_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@17 N_B[3]_XIbf3/MM1@17_d N_XIBF3/NET17_XIbf3/MM1@17_g
+ N_VSS_XIbf3/MM1@17_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@16 N_B[3]_XIbf3/MM1@16_d N_XIBF3/NET17_XIbf3/MM1@16_g
+ N_VSS_XIbf3/MM1@16_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@15 N_B[3]_XIbf3/MM1@15_d N_XIBF3/NET17_XIbf3/MM1@15_g
+ N_VSS_XIbf3/MM1@15_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@14 N_B[3]_XIbf3/MM1@14_d N_XIBF3/NET17_XIbf3/MM1@14_g
+ N_VSS_XIbf3/MM1@14_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@13 N_B[3]_XIbf3/MM1@13_d N_XIBF3/NET17_XIbf3/MM1@13_g
+ N_VSS_XIbf3/MM1@13_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@12 N_B[3]_XIbf3/MM1@12_d N_XIBF3/NET17_XIbf3/MM1@12_g
+ N_VSS_XIbf3/MM1@12_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@11 N_B[3]_XIbf3/MM1@11_d N_XIBF3/NET17_XIbf3/MM1@11_g
+ N_VSS_XIbf3/MM1@11_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@10 N_B[3]_XIbf3/MM1@10_d N_XIBF3/NET17_XIbf3/MM1@10_g
+ N_VSS_XIbf3/MM1@10_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@9 N_B[3]_XIbf3/MM1@9_d N_XIBF3/NET17_XIbf3/MM1@9_g
+ N_VSS_XIbf3/MM1@9_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@8 N_B[3]_XIbf3/MM1@8_d N_XIBF3/NET17_XIbf3/MM1@8_g
+ N_VSS_XIbf3/MM1@8_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@7 N_B[3]_XIbf3/MM1@7_d N_XIBF3/NET17_XIbf3/MM1@7_g
+ N_VSS_XIbf3/MM1@7_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@6 N_B[3]_XIbf3/MM1@6_d N_XIBF3/NET17_XIbf3/MM1@6_g
+ N_VSS_XIbf3/MM1@6_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@5 N_B[3]_XIbf3/MM1@5_d N_XIBF3/NET17_XIbf3/MM1@5_g
+ N_VSS_XIbf3/MM1@5_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@4 N_B[3]_XIbf3/MM1@4_d N_XIBF3/NET17_XIbf3/MM1@4_g
+ N_VSS_XIbf3/MM1@4_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@3 N_B[3]_XIbf3/MM1@3_d N_XIBF3/NET17_XIbf3/MM1@3_g
+ N_VSS_XIbf3/MM1@3_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM1@2 N_B[3]_XIbf3/MM1@2_d N_XIBF3/NET17_XIbf3/MM1@2_g
+ N_VSS_XIbf3/MM1@2_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mXIbf3/MM0 N_XIBF3/NET17_XIbf3/MM0_d N_NETB31_XIbf3/MM0_g N_VSS_XIbf3/MM0_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=7.35e-13 AS=3.825e-13 PD=2.48e-06
+ PS=5.1e-07
mXIbf3/MM0@7 N_XIBF3/NET17_XIbf3/MM0@7_d N_NETB31_XIbf3/MM0@7_g
+ N_VSS_XIbf3/MM0@7_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM0@6 N_XIBF3/NET17_XIbf3/MM0@6_d N_NETB31_XIbf3/MM0@6_g
+ N_VSS_XIbf3/MM0@6_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM0@5 N_XIBF3/NET17_XIbf3/MM0@5_d N_NETB31_XIbf3/MM0@5_g
+ N_VSS_XIbf3/MM0@5_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM0@4 N_XIBF3/NET17_XIbf3/MM0@4_d N_NETB31_XIbf3/MM0@4_g
+ N_VSS_XIbf3/MM0@4_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM0@3 N_XIBF3/NET17_XIbf3/MM0@3_d N_NETB31_XIbf3/MM0@3_g
+ N_VSS_XIbf3/MM0@3_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=3.825e-13 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM0@2 N_XIBF3/NET17_XIbf3/MM0@2_d N_NETB31_XIbf3/MM0@2_g
+ N_VSS_XIbf3/MM0@2_s N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=1.5e-06 AD=3.825e-13
+ AS=7.35e-13 PD=5.1e-07 PS=2.48e-06
mXI14/Mm2 N_INV14_XI14/Mm2_d N_T[14]_XI14/Mm2_g N_VSS_XI14/Mm2_s
+ N_VSS_XI01/MM1_b N_18 L=1.8e-07 W=2.08e-06 AD=1.0192e-12 AS=1.0192e-12
+ PD=3.06e-06 PS=3.06e-06
mXI01/MM2 N_ND01_XI01/MM2_d N_T[0]_XI01/MM2_g N_VDD_XI01/MM2_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXInd4/MM7 N_NETB1_XInd4/MM7_d N_ND13_XInd4/MM7_g N_VDD_XInd4/MM7_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=1.161e-05 AD=2.96055e-12 AS=5.6889e-12
+ PD=5.1e-07 PS=1.259e-05
mXI01/MM3 N_ND01_XI01/MM3_d N_INV1_XI01/MM3_g N_VDD_XI01/MM3_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXInd4/MM6 N_NETB1_XInd4/MM6_d N_ND57_XInd4/MM6_g N_VDD_XInd4/MM6_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=1.161e-05 AD=2.96055e-12 AS=2.96055e-12
+ PD=5.1e-07 PS=5.1e-07
mXInd4/MM5 N_NETB1_XInd4/MM5_d N_ND911_XInd4/MM5_g N_VDD_XInd4/MM5_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=1.161e-05 AD=2.96055e-12 AS=2.96055e-12
+ PD=5.1e-07 PS=5.1e-07
mXInd4/MM4 N_NETB1_XInd4/MM4_d N_INV13_XInd4/MM4_g N_VDD_XInd4/MM4_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=1.161e-05 AD=2.96055e-12 AS=5.6889e-12
+ PD=5.1e-07 PS=1.259e-05
mXI1/Mm1 N_INV1_XI1/Mm1_d N_T[1]_XI1/Mm1_g N_VDD_XI1/Mm1_s N_VDD_XI01/MM2_b P_18
+ L=1.8e-07 W=6.24e-06 AD=3.0576e-12 AS=3.0576e-12 PD=7.22e-06 PS=7.22e-06
mXInd22/MM3 N_NETB2_XInd22/MM3_d N_ND37_XInd22/MM3_g N_VDD_XInd22/MM3_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=1.625e-05 AD=4.14375e-12 AS=7.9625e-12
+ PD=5.1e-07 PS=1.723e-05
mXInd22/MM2 N_NETB2_XInd22/MM2_d N_INV11_XInd22/MM2_g N_VDD_XInd22/MM2_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=1.625e-05 AD=4.14375e-12 AS=7.9625e-12
+ PD=5.1e-07 PS=1.723e-05
mXInd13/MM2 N_ND13_XInd13/MM2_d N_T[1]_XInd13/MM2_g N_VDD_XInd13/MM2_s
+ N_VDD_XI01/MM2_b P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07
+ PS=5.98e-06
mXInd13/MM3 N_ND13_XInd13/MM3_d N_INV3_XInd13/MM3_g N_VDD_XInd13/MM3_s
+ N_VDD_XI01/MM2_b P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07
+ PS=5.98e-06
mXInd8/MM15 N_NETB0_XInd8/MM15_d N_INV14_XInd8/MM15_g N_VDD_XInd8/MM15_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=7.39e-06 AD=1.88445e-12 AS=3.6211e-12
+ PD=5.1e-07 PS=8.37e-06
mXInd8/MM14 N_NETB0_XInd8/MM14_d N_ND67_XInd8/MM14_g N_VDD_XInd8/MM14_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=7.39e-06 AD=1.88445e-12 AS=1.88445e-12
+ PD=5.1e-07 PS=5.1e-07
mXI23/MM2 N_ND23_XI23/MM2_d N_T[2]_XI23/MM2_g N_VDD_XI23/MM2_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXInd8/MM13 N_NETB0_XInd8/MM13_d N_ND01_XInd8/MM13_g N_VDD_XInd8/MM13_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=7.39e-06 AD=1.88445e-12 AS=1.88445e-12
+ PD=5.1e-07 PS=5.1e-07
mXI23/MM3 N_ND23_XI23/MM3_d N_INV3_XI23/MM3_g N_VDD_XI23/MM3_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXInd8/MM12 N_NETB0_XInd8/MM12_d N_ND23_XInd8/MM12_g N_VDD_XInd8/MM12_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=7.39e-06 AD=1.88445e-12 AS=1.88445e-12
+ PD=5.1e-07 PS=5.1e-07
mXInd8/MM11 N_NETB0_XInd8/MM11_d N_ND45_XInd8/MM11_g N_VDD_XInd8/MM11_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=7.39e-06 AD=1.88445e-12 AS=1.88445e-12
+ PD=5.1e-07 PS=5.1e-07
mXInd8/MM10 N_NETB0_XInd8/MM10_d N_ND89_XInd8/MM10_g N_VDD_XInd8/MM10_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=7.39e-06 AD=1.88445e-12 AS=1.88445e-12
+ PD=5.1e-07 PS=5.1e-07
mXI3/Mm1 N_INV3_XI3/Mm1_d N_T[3]_XI3/Mm1_g N_VDD_XI3/Mm1_s N_VDD_XI01/MM2_b P_18
+ L=1.8e-07 W=6.24e-06 AD=3.0576e-12 AS=3.0576e-12 PD=7.22e-06 PS=7.22e-06
mXInd8/MM8 N_NETB0_XInd8/MM8_d N_ND1011_XInd8/MM8_g N_VDD_XInd8/MM8_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=7.39e-06 AD=1.88445e-12 AS=1.88445e-12
+ PD=5.1e-07 PS=5.1e-07
mXInd8/MM9 N_NETB0_XInd8/MM9_d N_ND1213_XInd8/MM9_g N_VDD_XInd8/MM9_s
+ N_VDD_XInd4/MM7_b P_18 L=1.8e-07 W=7.39e-06 AD=1.88445e-12 AS=3.6211e-12
+ PD=5.1e-07 PS=8.37e-06
mXI37/MM2 N_ND37_XI37/MM2_d N_T[3]_XI37/MM2_g N_VDD_XI37/MM2_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXI37/MM3 N_ND37_XI37/MM3_d N_INV7_XI37/MM3_g N_VDD_XI37/MM3_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXI67/MM2 N_ND67_XI67/MM2_d N_T[6]_XI67/MM2_g N_VDD_XI67/MM2_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXI67/MM3 N_ND67_XI67/MM3_d N_INV7_XI67/MM3_g N_VDD_XI67/MM3_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXIbf0/MM3 N_B[0]_XIbf0/MM3_d N_XIBF0/NET17_XIbf0/MM3_g N_VDD_XIbf0/MM3_s
+ N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12 AS=2.205e-12
+ PD=5.1e-07 PS=5.48e-06
mXIbf0/MM3@28 N_B[0]_XIbf0/MM3@28_d N_XIBF0/NET17_XIbf0/MM3@28_g
+ N_VDD_XIbf0/MM3@28_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@27 N_B[0]_XIbf0/MM3@27_d N_XIBF0/NET17_XIbf0/MM3@27_g
+ N_VDD_XIbf0/MM3@27_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@26 N_B[0]_XIbf0/MM3@26_d N_XIBF0/NET17_XIbf0/MM3@26_g
+ N_VDD_XIbf0/MM3@26_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@25 N_B[0]_XIbf0/MM3@25_d N_XIBF0/NET17_XIbf0/MM3@25_g
+ N_VDD_XIbf0/MM3@25_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@24 N_B[0]_XIbf0/MM3@24_d N_XIBF0/NET17_XIbf0/MM3@24_g
+ N_VDD_XIbf0/MM3@24_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@23 N_B[0]_XIbf0/MM3@23_d N_XIBF0/NET17_XIbf0/MM3@23_g
+ N_VDD_XIbf0/MM3@23_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@22 N_B[0]_XIbf0/MM3@22_d N_XIBF0/NET17_XIbf0/MM3@22_g
+ N_VDD_XIbf0/MM3@22_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@21 N_B[0]_XIbf0/MM3@21_d N_XIBF0/NET17_XIbf0/MM3@21_g
+ N_VDD_XIbf0/MM3@21_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@20 N_B[0]_XIbf0/MM3@20_d N_XIBF0/NET17_XIbf0/MM3@20_g
+ N_VDD_XIbf0/MM3@20_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@19 N_B[0]_XIbf0/MM3@19_d N_XIBF0/NET17_XIbf0/MM3@19_g
+ N_VDD_XIbf0/MM3@19_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@18 N_B[0]_XIbf0/MM3@18_d N_XIBF0/NET17_XIbf0/MM3@18_g
+ N_VDD_XIbf0/MM3@18_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@17 N_B[0]_XIbf0/MM3@17_d N_XIBF0/NET17_XIbf0/MM3@17_g
+ N_VDD_XIbf0/MM3@17_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@16 N_B[0]_XIbf0/MM3@16_d N_XIBF0/NET17_XIbf0/MM3@16_g
+ N_VDD_XIbf0/MM3@16_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@15 N_B[0]_XIbf0/MM3@15_d N_XIBF0/NET17_XIbf0/MM3@15_g
+ N_VDD_XIbf0/MM3@15_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@14 N_B[0]_XIbf0/MM3@14_d N_XIBF0/NET17_XIbf0/MM3@14_g
+ N_VDD_XIbf0/MM3@14_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@13 N_B[0]_XIbf0/MM3@13_d N_XIBF0/NET17_XIbf0/MM3@13_g
+ N_VDD_XIbf0/MM3@13_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@12 N_B[0]_XIbf0/MM3@12_d N_XIBF0/NET17_XIbf0/MM3@12_g
+ N_VDD_XIbf0/MM3@12_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@11 N_B[0]_XIbf0/MM3@11_d N_XIBF0/NET17_XIbf0/MM3@11_g
+ N_VDD_XIbf0/MM3@11_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@10 N_B[0]_XIbf0/MM3@10_d N_XIBF0/NET17_XIbf0/MM3@10_g
+ N_VDD_XIbf0/MM3@10_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@9 N_B[0]_XIbf0/MM3@9_d N_XIBF0/NET17_XIbf0/MM3@9_g
+ N_VDD_XIbf0/MM3@9_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@8 N_B[0]_XIbf0/MM3@8_d N_XIBF0/NET17_XIbf0/MM3@8_g
+ N_VDD_XIbf0/MM3@8_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@7 N_B[0]_XIbf0/MM3@7_d N_XIBF0/NET17_XIbf0/MM3@7_g
+ N_VDD_XIbf0/MM3@7_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@6 N_B[0]_XIbf0/MM3@6_d N_XIBF0/NET17_XIbf0/MM3@6_g
+ N_VDD_XIbf0/MM3@6_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@5 N_B[0]_XIbf0/MM3@5_d N_XIBF0/NET17_XIbf0/MM3@5_g
+ N_VDD_XIbf0/MM3@5_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@4 N_B[0]_XIbf0/MM3@4_d N_XIBF0/NET17_XIbf0/MM3@4_g
+ N_VDD_XIbf0/MM3@4_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@3 N_B[0]_XIbf0/MM3@3_d N_XIBF0/NET17_XIbf0/MM3@3_g
+ N_VDD_XIbf0/MM3@3_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM3@2 N_B[0]_XIbf0/MM3@2_d N_XIBF0/NET17_XIbf0/MM3@2_g
+ N_VDD_XIbf0/MM3@2_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=2.205e-12 PD=5.1e-07 PS=5.48e-06
mXIbf0/MM2 N_XIBF0/NET17_XIbf0/MM2_d N_NETB0_XIbf0/MM2_g N_VDD_XIbf0/MM2_s
+ N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=2.205e-12 AS=1.1475e-12
+ PD=5.48e-06 PS=5.1e-07
mXIbf0/MM2@7 N_XIBF0/NET17_XIbf0/MM2@7_d N_NETB0_XIbf0/MM2@7_g
+ N_VDD_XIbf0/MM2@7_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM2@6 N_XIBF0/NET17_XIbf0/MM2@6_d N_NETB0_XIbf0/MM2@6_g
+ N_VDD_XIbf0/MM2@6_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM2@5 N_XIBF0/NET17_XIbf0/MM2@5_d N_NETB0_XIbf0/MM2@5_g
+ N_VDD_XIbf0/MM2@5_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM2@4 N_XIBF0/NET17_XIbf0/MM2@4_d N_NETB0_XIbf0/MM2@4_g
+ N_VDD_XIbf0/MM2@4_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM2@3 N_XIBF0/NET17_XIbf0/MM2@3_d N_NETB0_XIbf0/MM2@3_g
+ N_VDD_XIbf0/MM2@3_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf0/MM2@2 N_XIBF0/NET17_XIbf0/MM2@2_d N_NETB0_XIbf0/MM2@2_g
+ N_VDD_XIbf0/MM2@2_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=2.205e-12 PD=5.1e-07 PS=5.48e-06
mXIb31/Mm1 N_NETB31_XIb31/Mm1_d N_INV7_XIb31/Mm1_g N_VDD_XIb31/Mm1_s
+ N_VDD_XI01/MM2_b P_18 L=1.8e-07 W=6.24e-06 AD=3.0576e-12 AS=3.0576e-12
+ PD=7.22e-06 PS=7.22e-06
mXI7/Mm1 N_INV7_XI7/Mm1_d N_T[7]_XI7/Mm1_g N_VDD_XI7/Mm1_s N_VDD_XI01/MM2_b P_18
+ L=1.8e-07 W=6.24e-06 AD=3.0576e-12 AS=3.0576e-12 PD=7.22e-06 PS=7.22e-06
mXI57/MM3 N_ND57_XI57/MM3_d N_INV7_XI57/MM3_g N_VDD_XI57/MM3_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXIbf1/MM3 N_B[1]_XIbf1/MM3_d N_XIBF1/NET17_XIbf1/MM3_g N_VDD_XIbf1/MM3_s
+ N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12 AS=2.205e-12
+ PD=5.1e-07 PS=5.48e-06
mXIbf1/MM3@28 N_B[1]_XIbf1/MM3@28_d N_XIBF1/NET17_XIbf1/MM3@28_g
+ N_VDD_XIbf1/MM3@28_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@27 N_B[1]_XIbf1/MM3@27_d N_XIBF1/NET17_XIbf1/MM3@27_g
+ N_VDD_XIbf1/MM3@27_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@26 N_B[1]_XIbf1/MM3@26_d N_XIBF1/NET17_XIbf1/MM3@26_g
+ N_VDD_XIbf1/MM3@26_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@25 N_B[1]_XIbf1/MM3@25_d N_XIBF1/NET17_XIbf1/MM3@25_g
+ N_VDD_XIbf1/MM3@25_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@24 N_B[1]_XIbf1/MM3@24_d N_XIBF1/NET17_XIbf1/MM3@24_g
+ N_VDD_XIbf1/MM3@24_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@23 N_B[1]_XIbf1/MM3@23_d N_XIBF1/NET17_XIbf1/MM3@23_g
+ N_VDD_XIbf1/MM3@23_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@22 N_B[1]_XIbf1/MM3@22_d N_XIBF1/NET17_XIbf1/MM3@22_g
+ N_VDD_XIbf1/MM3@22_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@21 N_B[1]_XIbf1/MM3@21_d N_XIBF1/NET17_XIbf1/MM3@21_g
+ N_VDD_XIbf1/MM3@21_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@20 N_B[1]_XIbf1/MM3@20_d N_XIBF1/NET17_XIbf1/MM3@20_g
+ N_VDD_XIbf1/MM3@20_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@19 N_B[1]_XIbf1/MM3@19_d N_XIBF1/NET17_XIbf1/MM3@19_g
+ N_VDD_XIbf1/MM3@19_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@18 N_B[1]_XIbf1/MM3@18_d N_XIBF1/NET17_XIbf1/MM3@18_g
+ N_VDD_XIbf1/MM3@18_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@17 N_B[1]_XIbf1/MM3@17_d N_XIBF1/NET17_XIbf1/MM3@17_g
+ N_VDD_XIbf1/MM3@17_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@16 N_B[1]_XIbf1/MM3@16_d N_XIBF1/NET17_XIbf1/MM3@16_g
+ N_VDD_XIbf1/MM3@16_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@15 N_B[1]_XIbf1/MM3@15_d N_XIBF1/NET17_XIbf1/MM3@15_g
+ N_VDD_XIbf1/MM3@15_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@14 N_B[1]_XIbf1/MM3@14_d N_XIBF1/NET17_XIbf1/MM3@14_g
+ N_VDD_XIbf1/MM3@14_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@13 N_B[1]_XIbf1/MM3@13_d N_XIBF1/NET17_XIbf1/MM3@13_g
+ N_VDD_XIbf1/MM3@13_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@12 N_B[1]_XIbf1/MM3@12_d N_XIBF1/NET17_XIbf1/MM3@12_g
+ N_VDD_XIbf1/MM3@12_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@11 N_B[1]_XIbf1/MM3@11_d N_XIBF1/NET17_XIbf1/MM3@11_g
+ N_VDD_XIbf1/MM3@11_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@10 N_B[1]_XIbf1/MM3@10_d N_XIBF1/NET17_XIbf1/MM3@10_g
+ N_VDD_XIbf1/MM3@10_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@9 N_B[1]_XIbf1/MM3@9_d N_XIBF1/NET17_XIbf1/MM3@9_g
+ N_VDD_XIbf1/MM3@9_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@8 N_B[1]_XIbf1/MM3@8_d N_XIBF1/NET17_XIbf1/MM3@8_g
+ N_VDD_XIbf1/MM3@8_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@7 N_B[1]_XIbf1/MM3@7_d N_XIBF1/NET17_XIbf1/MM3@7_g
+ N_VDD_XIbf1/MM3@7_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@6 N_B[1]_XIbf1/MM3@6_d N_XIBF1/NET17_XIbf1/MM3@6_g
+ N_VDD_XIbf1/MM3@6_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@5 N_B[1]_XIbf1/MM3@5_d N_XIBF1/NET17_XIbf1/MM3@5_g
+ N_VDD_XIbf1/MM3@5_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@4 N_B[1]_XIbf1/MM3@4_d N_XIBF1/NET17_XIbf1/MM3@4_g
+ N_VDD_XIbf1/MM3@4_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@3 N_B[1]_XIbf1/MM3@3_d N_XIBF1/NET17_XIbf1/MM3@3_g
+ N_VDD_XIbf1/MM3@3_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM3@2 N_B[1]_XIbf1/MM3@2_d N_XIBF1/NET17_XIbf1/MM3@2_g
+ N_VDD_XIbf1/MM3@2_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=2.205e-12 PD=5.1e-07 PS=5.48e-06
mXIbf1/MM2 N_XIBF1/NET17_XIbf1/MM2_d N_NETB1_XIbf1/MM2_g N_VDD_XIbf1/MM2_s
+ N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=2.205e-12 AS=1.1475e-12
+ PD=5.48e-06 PS=5.1e-07
mXIbf1/MM2@7 N_XIBF1/NET17_XIbf1/MM2@7_d N_NETB1_XIbf1/MM2@7_g
+ N_VDD_XIbf1/MM2@7_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM2@6 N_XIBF1/NET17_XIbf1/MM2@6_d N_NETB1_XIbf1/MM2@6_g
+ N_VDD_XIbf1/MM2@6_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM2@5 N_XIBF1/NET17_XIbf1/MM2@5_d N_NETB1_XIbf1/MM2@5_g
+ N_VDD_XIbf1/MM2@5_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM2@4 N_XIBF1/NET17_XIbf1/MM2@4_d N_NETB1_XIbf1/MM2@4_g
+ N_VDD_XIbf1/MM2@4_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM2@3 N_XIBF1/NET17_XIbf1/MM2@3_d N_NETB1_XIbf1/MM2@3_g
+ N_VDD_XIbf1/MM2@3_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf1/MM2@2 N_XIBF1/NET17_XIbf1/MM2@2_d N_NETB1_XIbf1/MM2@2_g
+ N_VDD_XIbf1/MM2@2_s N_VDD_XIbf0/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=2.205e-12 PD=5.1e-07 PS=5.48e-06
mXI57/MM2 N_ND57_XI57/MM2_d N_T[5]_XI57/MM2_g N_VDD_XI57/MM2_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXI5/Mm1 N_INV5_XI5/Mm1_d N_T[5]_XI5/Mm1_g N_VDD_XI5/Mm1_s N_VDD_XI01/MM2_b P_18
+ L=1.8e-07 W=6.24e-06 AD=3.0576e-12 AS=3.0576e-12 PD=7.22e-06 PS=7.22e-06
mXI45/MM3 N_ND45_XI45/MM3_d N_INV5_XI45/MM3_g N_VDD_XI45/MM3_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXI45/MM2 N_ND45_XI45/MM2_d N_T[4]_XI45/MM2_g N_VDD_XI45/MM2_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXI89/MM2 N_ND89_XI89/MM2_d N_T[8]_XI89/MM2_g N_VDD_XI89/MM2_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXI89/MM3 N_ND89_XI89/MM3_d N_INV9_XI89/MM3_g N_VDD_XI89/MM3_s N_VDD_XI01/MM2_b
+ P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07 PS=5.98e-06
mXI9/Mm1 N_INV9_XI9/Mm1_d N_T[9]_XI9/Mm1_g N_VDD_XI9/Mm1_s N_VDD_XI01/MM2_b P_18
+ L=1.8e-07 W=6.24e-06 AD=3.0576e-12 AS=3.0576e-12 PD=7.22e-06 PS=7.22e-06
mXIbf2/MM3 N_B[2]_XIbf2/MM3_d N_XIBF2/NET17_XIbf2/MM3_g N_VDD_XIbf2/MM3_s
+ N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12 AS=2.205e-12
+ PD=5.1e-07 PS=5.48e-06
mXIbf2/MM3@28 N_B[2]_XIbf2/MM3@28_d N_XIBF2/NET17_XIbf2/MM3@28_g
+ N_VDD_XIbf2/MM3@28_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@27 N_B[2]_XIbf2/MM3@27_d N_XIBF2/NET17_XIbf2/MM3@27_g
+ N_VDD_XIbf2/MM3@27_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@26 N_B[2]_XIbf2/MM3@26_d N_XIBF2/NET17_XIbf2/MM3@26_g
+ N_VDD_XIbf2/MM3@26_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@25 N_B[2]_XIbf2/MM3@25_d N_XIBF2/NET17_XIbf2/MM3@25_g
+ N_VDD_XIbf2/MM3@25_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@24 N_B[2]_XIbf2/MM3@24_d N_XIBF2/NET17_XIbf2/MM3@24_g
+ N_VDD_XIbf2/MM3@24_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@23 N_B[2]_XIbf2/MM3@23_d N_XIBF2/NET17_XIbf2/MM3@23_g
+ N_VDD_XIbf2/MM3@23_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@22 N_B[2]_XIbf2/MM3@22_d N_XIBF2/NET17_XIbf2/MM3@22_g
+ N_VDD_XIbf2/MM3@22_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@21 N_B[2]_XIbf2/MM3@21_d N_XIBF2/NET17_XIbf2/MM3@21_g
+ N_VDD_XIbf2/MM3@21_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@20 N_B[2]_XIbf2/MM3@20_d N_XIBF2/NET17_XIbf2/MM3@20_g
+ N_VDD_XIbf2/MM3@20_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@19 N_B[2]_XIbf2/MM3@19_d N_XIBF2/NET17_XIbf2/MM3@19_g
+ N_VDD_XIbf2/MM3@19_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@18 N_B[2]_XIbf2/MM3@18_d N_XIBF2/NET17_XIbf2/MM3@18_g
+ N_VDD_XIbf2/MM3@18_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@17 N_B[2]_XIbf2/MM3@17_d N_XIBF2/NET17_XIbf2/MM3@17_g
+ N_VDD_XIbf2/MM3@17_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@16 N_B[2]_XIbf2/MM3@16_d N_XIBF2/NET17_XIbf2/MM3@16_g
+ N_VDD_XIbf2/MM3@16_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@15 N_B[2]_XIbf2/MM3@15_d N_XIBF2/NET17_XIbf2/MM3@15_g
+ N_VDD_XIbf2/MM3@15_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@14 N_B[2]_XIbf2/MM3@14_d N_XIBF2/NET17_XIbf2/MM3@14_g
+ N_VDD_XIbf2/MM3@14_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@13 N_B[2]_XIbf2/MM3@13_d N_XIBF2/NET17_XIbf2/MM3@13_g
+ N_VDD_XIbf2/MM3@13_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@12 N_B[2]_XIbf2/MM3@12_d N_XIBF2/NET17_XIbf2/MM3@12_g
+ N_VDD_XIbf2/MM3@12_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@11 N_B[2]_XIbf2/MM3@11_d N_XIBF2/NET17_XIbf2/MM3@11_g
+ N_VDD_XIbf2/MM3@11_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@10 N_B[2]_XIbf2/MM3@10_d N_XIBF2/NET17_XIbf2/MM3@10_g
+ N_VDD_XIbf2/MM3@10_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@9 N_B[2]_XIbf2/MM3@9_d N_XIBF2/NET17_XIbf2/MM3@9_g
+ N_VDD_XIbf2/MM3@9_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@8 N_B[2]_XIbf2/MM3@8_d N_XIBF2/NET17_XIbf2/MM3@8_g
+ N_VDD_XIbf2/MM3@8_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@7 N_B[2]_XIbf2/MM3@7_d N_XIBF2/NET17_XIbf2/MM3@7_g
+ N_VDD_XIbf2/MM3@7_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@6 N_B[2]_XIbf2/MM3@6_d N_XIBF2/NET17_XIbf2/MM3@6_g
+ N_VDD_XIbf2/MM3@6_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@5 N_B[2]_XIbf2/MM3@5_d N_XIBF2/NET17_XIbf2/MM3@5_g
+ N_VDD_XIbf2/MM3@5_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@4 N_B[2]_XIbf2/MM3@4_d N_XIBF2/NET17_XIbf2/MM3@4_g
+ N_VDD_XIbf2/MM3@4_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@3 N_B[2]_XIbf2/MM3@3_d N_XIBF2/NET17_XIbf2/MM3@3_g
+ N_VDD_XIbf2/MM3@3_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM3@2 N_B[2]_XIbf2/MM3@2_d N_XIBF2/NET17_XIbf2/MM3@2_g
+ N_VDD_XIbf2/MM3@2_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=2.205e-12 PD=5.1e-07 PS=5.48e-06
mXIbf2/MM2 N_XIBF2/NET17_XIbf2/MM2_d N_NETB2_XIbf2/MM2_g N_VDD_XIbf2/MM2_s
+ N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=2.205e-12 AS=1.1475e-12
+ PD=5.48e-06 PS=5.1e-07
mXIbf2/MM2@7 N_XIBF2/NET17_XIbf2/MM2@7_d N_NETB2_XIbf2/MM2@7_g
+ N_VDD_XIbf2/MM2@7_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM2@6 N_XIBF2/NET17_XIbf2/MM2@6_d N_NETB2_XIbf2/MM2@6_g
+ N_VDD_XIbf2/MM2@6_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM2@5 N_XIBF2/NET17_XIbf2/MM2@5_d N_NETB2_XIbf2/MM2@5_g
+ N_VDD_XIbf2/MM2@5_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM2@4 N_XIBF2/NET17_XIbf2/MM2@4_d N_NETB2_XIbf2/MM2@4_g
+ N_VDD_XIbf2/MM2@4_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM2@3 N_XIBF2/NET17_XIbf2/MM2@3_d N_NETB2_XIbf2/MM2@3_g
+ N_VDD_XIbf2/MM2@3_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf2/MM2@2 N_XIBF2/NET17_XIbf2/MM2@2_d N_NETB2_XIbf2/MM2@2_g
+ N_VDD_XIbf2/MM2@2_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=2.205e-12 PD=5.1e-07 PS=5.48e-06
mXI911/MM2 N_ND911_XI911/MM2_d N_T[9]_XI911/MM2_g N_VDD_XI911/MM2_s
+ N_VDD_XI01/MM2_b P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07
+ PS=5.98e-06
mXI911/MM3 N_ND911_XI911/MM3_d N_INV11_XI911/MM3_g N_VDD_XI911/MM3_s
+ N_VDD_XI01/MM2_b P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07
+ PS=5.98e-06
mXI1011/MM2 N_ND1011_XI1011/MM2_d N_T[10]_XI1011/MM2_g N_VDD_XI1011/MM2_s
+ N_VDD_XI01/MM2_b P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07
+ PS=5.98e-06
mXI1011/MM3 N_ND1011_XI1011/MM3_d N_INV11_XI1011/MM3_g N_VDD_XI1011/MM3_s
+ N_VDD_XI01/MM2_b P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07
+ PS=5.98e-06
mXI11/Mm1 N_INV11_XI11/Mm1_d N_T[11]_XI11/Mm1_g N_VDD_XI11/Mm1_s
+ N_VDD_XI01/MM2_b P_18 L=1.8e-07 W=6.24e-06 AD=3.0576e-12 AS=3.0576e-12
+ PD=7.22e-06 PS=7.22e-06
mXIbf3/MM3 N_B[3]_XIbf3/MM3_d N_XIBF3/NET17_XIbf3/MM3_g N_VDD_XIbf3/MM3_s
+ N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12 AS=2.205e-12
+ PD=5.1e-07 PS=5.48e-06
mXIbf3/MM3@28 N_B[3]_XIbf3/MM3@28_d N_XIBF3/NET17_XIbf3/MM3@28_g
+ N_VDD_XIbf3/MM3@28_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@27 N_B[3]_XIbf3/MM3@27_d N_XIBF3/NET17_XIbf3/MM3@27_g
+ N_VDD_XIbf3/MM3@27_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@26 N_B[3]_XIbf3/MM3@26_d N_XIBF3/NET17_XIbf3/MM3@26_g
+ N_VDD_XIbf3/MM3@26_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@25 N_B[3]_XIbf3/MM3@25_d N_XIBF3/NET17_XIbf3/MM3@25_g
+ N_VDD_XIbf3/MM3@25_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@24 N_B[3]_XIbf3/MM3@24_d N_XIBF3/NET17_XIbf3/MM3@24_g
+ N_VDD_XIbf3/MM3@24_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@23 N_B[3]_XIbf3/MM3@23_d N_XIBF3/NET17_XIbf3/MM3@23_g
+ N_VDD_XIbf3/MM3@23_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@22 N_B[3]_XIbf3/MM3@22_d N_XIBF3/NET17_XIbf3/MM3@22_g
+ N_VDD_XIbf3/MM3@22_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@21 N_B[3]_XIbf3/MM3@21_d N_XIBF3/NET17_XIbf3/MM3@21_g
+ N_VDD_XIbf3/MM3@21_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@20 N_B[3]_XIbf3/MM3@20_d N_XIBF3/NET17_XIbf3/MM3@20_g
+ N_VDD_XIbf3/MM3@20_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@19 N_B[3]_XIbf3/MM3@19_d N_XIBF3/NET17_XIbf3/MM3@19_g
+ N_VDD_XIbf3/MM3@19_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@18 N_B[3]_XIbf3/MM3@18_d N_XIBF3/NET17_XIbf3/MM3@18_g
+ N_VDD_XIbf3/MM3@18_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@17 N_B[3]_XIbf3/MM3@17_d N_XIBF3/NET17_XIbf3/MM3@17_g
+ N_VDD_XIbf3/MM3@17_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@16 N_B[3]_XIbf3/MM3@16_d N_XIBF3/NET17_XIbf3/MM3@16_g
+ N_VDD_XIbf3/MM3@16_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@15 N_B[3]_XIbf3/MM3@15_d N_XIBF3/NET17_XIbf3/MM3@15_g
+ N_VDD_XIbf3/MM3@15_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@14 N_B[3]_XIbf3/MM3@14_d N_XIBF3/NET17_XIbf3/MM3@14_g
+ N_VDD_XIbf3/MM3@14_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@13 N_B[3]_XIbf3/MM3@13_d N_XIBF3/NET17_XIbf3/MM3@13_g
+ N_VDD_XIbf3/MM3@13_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@12 N_B[3]_XIbf3/MM3@12_d N_XIBF3/NET17_XIbf3/MM3@12_g
+ N_VDD_XIbf3/MM3@12_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@11 N_B[3]_XIbf3/MM3@11_d N_XIBF3/NET17_XIbf3/MM3@11_g
+ N_VDD_XIbf3/MM3@11_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@10 N_B[3]_XIbf3/MM3@10_d N_XIBF3/NET17_XIbf3/MM3@10_g
+ N_VDD_XIbf3/MM3@10_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@9 N_B[3]_XIbf3/MM3@9_d N_XIBF3/NET17_XIbf3/MM3@9_g
+ N_VDD_XIbf3/MM3@9_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@8 N_B[3]_XIbf3/MM3@8_d N_XIBF3/NET17_XIbf3/MM3@8_g
+ N_VDD_XIbf3/MM3@8_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@7 N_B[3]_XIbf3/MM3@7_d N_XIBF3/NET17_XIbf3/MM3@7_g
+ N_VDD_XIbf3/MM3@7_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@6 N_B[3]_XIbf3/MM3@6_d N_XIBF3/NET17_XIbf3/MM3@6_g
+ N_VDD_XIbf3/MM3@6_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@5 N_B[3]_XIbf3/MM3@5_d N_XIBF3/NET17_XIbf3/MM3@5_g
+ N_VDD_XIbf3/MM3@5_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@4 N_B[3]_XIbf3/MM3@4_d N_XIBF3/NET17_XIbf3/MM3@4_g
+ N_VDD_XIbf3/MM3@4_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@3 N_B[3]_XIbf3/MM3@3_d N_XIBF3/NET17_XIbf3/MM3@3_g
+ N_VDD_XIbf3/MM3@3_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM3@2 N_B[3]_XIbf3/MM3@2_d N_XIBF3/NET17_XIbf3/MM3@2_g
+ N_VDD_XIbf3/MM3@2_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=2.205e-12 PD=5.1e-07 PS=5.48e-06
mXIbf3/MM2 N_XIBF3/NET17_XIbf3/MM2_d N_NETB31_XIbf3/MM2_g N_VDD_XIbf3/MM2_s
+ N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=2.205e-12 AS=1.1475e-12
+ PD=5.48e-06 PS=5.1e-07
mXIbf3/MM2@7 N_XIBF3/NET17_XIbf3/MM2@7_d N_NETB31_XIbf3/MM2@7_g
+ N_VDD_XIbf3/MM2@7_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM2@6 N_XIBF3/NET17_XIbf3/MM2@6_d N_NETB31_XIbf3/MM2@6_g
+ N_VDD_XIbf3/MM2@6_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM2@5 N_XIBF3/NET17_XIbf3/MM2@5_d N_NETB31_XIbf3/MM2@5_g
+ N_VDD_XIbf3/MM2@5_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM2@4 N_XIBF3/NET17_XIbf3/MM2@4_d N_NETB31_XIbf3/MM2@4_g
+ N_VDD_XIbf3/MM2@4_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM2@3 N_XIBF3/NET17_XIbf3/MM2@3_d N_NETB31_XIbf3/MM2@3_g
+ N_VDD_XIbf3/MM2@3_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=1.1475e-12 PD=5.1e-07 PS=5.1e-07
mXIbf3/MM2@2 N_XIBF3/NET17_XIbf3/MM2@2_d N_NETB31_XIbf3/MM2@2_g
+ N_VDD_XIbf3/MM2@2_s N_VDD_XIbf2/MM3_b P_18 L=1.8e-07 W=4.5e-06 AD=1.1475e-12
+ AS=2.205e-12 PD=5.1e-07 PS=5.48e-06
mXI1213/MM2 N_ND1213_XI1213/MM2_d N_T[12]_XI1213/MM2_g N_VDD_XI1213/MM2_s
+ N_VDD_XI01/MM2_b P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07
+ PS=5.98e-06
mXI1213/MM3 N_ND1213_XI1213/MM3_d N_INV13_XI1213/MM3_g N_VDD_XI1213/MM3_s
+ N_VDD_XI01/MM2_b P_18 L=1.8e-07 W=5e-06 AD=1.275e-12 AS=2.45e-12 PD=5.1e-07
+ PS=5.98e-06
mXI13/Mm1 N_INV13_XI13/Mm1_d N_T[13]_XI13/Mm1_g N_VDD_XI13/Mm1_s
+ N_VDD_XI01/MM2_b P_18 L=1.8e-07 W=6.24e-06 AD=3.0576e-12 AS=3.0576e-12
+ PD=7.22e-06 PS=7.22e-06
mXI14/Mm1 N_INV14_XI14/Mm1_d N_T[14]_XI14/Mm1_g N_VDD_XI14/Mm1_s
+ N_VDD_XI01/MM2_b P_18 L=1.8e-07 W=6.24e-06 AD=3.0576e-12 AS=3.0576e-12
+ PD=7.22e-06 PS=7.22e-06
*
.include "TBC.pex.spi.TBC.pxi"
*
.ends
*
*
