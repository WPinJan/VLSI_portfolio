************************************************************************
* auCdl Netlist:
* 
* Library Name:  VLSI
* Top Cell Name: TBC2
* View Name:     schematic
* Netlisted on:  Oct 24 22:04:44 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.param Ln= 0.18u
.param Lp= 0.18u


.param Wninv= 2.08u
.param Wpinv= 6.24u
.param Wnnand2= 3.32u
.param Wpnand2= 5.00u

.param Wnnand22= 10.84u
.param Wpnand22= 16.25u
.param Wnnand4= 15.48u
.param Wpnand4= 11.61u
.param Wnnand8= 19.70u
.param Wpnand8= 7.39u
.param WninvB01= 1.5u
.param WpinvB01= 4.5u
.param WninvB02= 1.5u
.param WpinvB02= 4.5u


************************************************************************
* Library Name: VLSI
* Cell Name:    NAND8
* View Name:    schematic
************************************************************************

.SUBCKT NAND8 A B C D E F G H OUT VDD VSS
*.PININFO A:I B:I C:I D:I E:I F:I G:I H:I OUT:O VDD:B VSS:B
MM15 OUT H VDD VDD P_18 W=Wpnand8 L=Lp m=1
MM14 OUT G VDD VDD P_18 W=Wpnand8 L=Lp m=1
MM13 OUT F VDD VDD P_18 W=Wpnand8 L=Lp m=1
MM12 OUT E VDD VDD P_18 W=Wpnand8 L=Lp m=1
MM11 OUT D VDD VDD P_18 W=Wpnand8 L=Lp m=1
MM10 OUT C VDD VDD P_18 W=Wpnand8 L=Lp m=1
MM9 OUT B VDD VDD P_18 W=Wpnand8 L=Lp m=1
MM8 OUT A VDD VDD P_18 W=Wpnand8 L=Lp m=1
MM7 net44 H VSS VSS N_18 W=Wnnand8 L=Ln m=1
MM6 net48 G net44 VSS N_18 W=Wnnand8 L=Ln m=1
MM5 net52 F net48 VSS N_18 W=Wnnand8 L=Ln m=1
MM4 net56 E net52 VSS N_18 W=Wnnand8 L=Ln m=1
MM3 net60 D net56 VSS N_18 W=Wnnand8 L=Ln m=1
MM2 net64 C net60 VSS N_18 W=Wnnand8 L=Ln m=1
MM1 net68 B net64 VSS N_18 W=Wnnand8 L=Ln m=1
MM0 OUT A net68 VSS N_18 W=Wnnand8 L=Ln m=1
.ENDS

************************************************************************
* Library Name: VLSI
* Cell Name:    NAND4
* View Name:    schematic
************************************************************************

.SUBCKT NAND4 A B C D OUT VDD VSS
*.PININFO A:I B:I C:I D:I OUT:O VDD:B VSS:B
MM7 OUT D VDD VDD P_18 W=Wpnand4 L=Lp m=1
MM6 OUT C VDD VDD P_18 W=Wpnand4 L=Lp m=1
MM5 OUT B VDD VDD P_18 W=Wpnand4 L=Lp m=1
MM4 OUT A VDD VDD P_18 W=Wpnand4 L=Lp m=1
MM3 net24 D VSS VSS N_18 W=Wnnand4 L=Ln m=1
MM2 net28 C net24 VSS N_18 W=Wnnand4 L=Ln m=1
MM1 net32 B net28 VSS N_18 W=Wnnand4 L=Ln m=1
MM0 OUT A net32 VSS N_18 W=Wnnand4 L=Ln m=1
.ENDS

************************************************************************
* Library Name: VLSI
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VOUT VSS
*.PININFO A:I B:I VOUT:O VDD:B VSS:B
MM2 VOUT B VDD VDD P_18 W=Wpnand2 L=Lp m=1
MM3 VOUT A VDD VDD P_18 W=Wpnand2 L=Lp m=1
MM0 VOUT A net14 VSS N_18 W=Wnnand2 L=Ln m=1
MM1 net14 B VSS VSS N_18 W=Wnnand2 L=Ln m=1
.ENDS

.SUBCKT NAND22 A B VDD VOUT VSS
*.PININFO A:I B:I VOUT:O VDD:B VSS:B
MM2 VOUT B VDD VDD P_18 W=Wpnand22 L=Lp m=1
MM3 VOUT A VDD VDD P_18 W=Wpnand22 L=Lp m=1
MM0 VOUT A net14 VSS N_18 W=Wnnand22 L=Ln m=1
MM1 net14 B VSS VSS N_18 W=Wnnand22 L=Ln m=1
.ENDS

************************************************************************
* Library Name: VLSI
* Cell Name:    inv
* View Name:    schematic
************************************************************************

.SUBCKT inv IN OUT VDD VSS
*.PININFO IN:I OUT:O VDD:B VSS:B
Mm2 OUT IN VSS VSS N_18 W=Wninv L=Ln m=1
Mm1 OUT IN VDD VDD P_18 W=Wpinv L=Lp m=1
.ENDS


************************************************************************
* Library Name: VLSI
* Cell Name:    buff
* View Name:    schematic
************************************************************************

.SUBCKT buffB0 VDD VSS in out
*.PININFO in:I out:O VDD:B VSS:B
MM3 out net17 VDD VDD P_18 W=WpinvB02 L=Lp m=28
MM2 net17 in VDD VDD P_18 W=WpinvB01 L=Lp m=7
MM1 out net17 VSS VSS N_18 W=WninvB02 L=Ln m=28
MM0 net17 in VSS VSS N_18 W=WninvB01 L=Ln m=7
.ENDS


************************************************************************
* Library Name: VLSI
* Cell Name:    TBC2
* View Name:    schematic
************************************************************************

.SUBCKT TBC VDD VSS T[0] T[1] T[2] T[3] T[4] T[5] T[6] T[7] T[8] T[9] T[10] T[11] T[12]
+ T[13] T[14] B[0] B[1] B[2] B[3]
*.PININFO T[0]:I T[1]:I T[2]:I T[3]:I T[4]:I T[5]:I T[6]:I T[7]:I T[8]:I 
*.PININFO T[9]:I T[10]:I T[11]:I T[12]:I T[13]:I T[14]:I B[0]:O B[1]:O B[2]:O 
*.PININFO B[3]:O VDD:B VSS:B


XI01 inv1 T[0] VDD nd01 VSS / NAND2
XI1 T[1] inv1 VDD VSS / inv
XInd13 inv3 T[1] VDD nd13 VSS / NAND2
XI23 inv3 T[2] VDD nd23 VSS / NAND2
XI3 T[3] inv3 VDD VSS / inv
XI37 inv7 T[3] VDD nd37 VSS / NAND2
XI45 inv5 T[4] VDD nd45 VSS / NAND2
XI5 T[5] inv5 VDD VSS / inv
XI57 inv7 T[5] VDD nd57 VSS / NAND2
XI67 inv7 T[6] VDD nd67 VSS / NAND2
XI7 T[7] inv7 VDD VSS / inv
XI89 inv9 T[8] VDD nd89 VSS / NAND2
XI9 T[9] inv9 VDD VSS / inv
XI911 inv11 T[9] VDD nd911 VSS / NAND2
XI1011 inv11 T[10] VDD nd1011 VSS / NAND2
XI11 T[11] inv11 VDD VSS / inv
XI1213 inv13 T[12] VDD nd1213 VSS / NAND2
XI13 T[13] inv13 VDD VSS / inv
XI14 T[14] inv14 VDD VSS / inv


XInd22 nd37 inv11 VDD netB2 VSS / NAND22
XInd4  inv13 nd911 nd57 nd13 netB1 VDD VSS / NAND4
XInd8  nd1213 nd1011 nd89 nd45 nd23 nd01 nd67 inv14 netB0 VDD VSS / 
+ NAND8
XIbf0 VDD VSS netB0 B[0] / buffB0
XIbf1 VDD VSS netB1 B[1] / buffB0
XIbf2 VDD VSS netB2 B[2] / buffB0
XIb31 inv7 netb31 VDD VSS / inv
XIbf3 VDD VSS netb31 B[3] / buffB0

.ENDS










