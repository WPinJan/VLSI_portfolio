************************************************************************
* auCdl Netlist:
* 
* Library Name:  VLSI
* Top Cell Name: DFFnand
* View Name:     schematic
* Netlisted on:  Nov 13 15:45:19 2024
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM


************************************************************************
* Library Name: VLSI
* Cell Name:    inv
* View Name:    schematic
************************************************************************

.SUBCKT inv IN OUT VDD VSS
*.PININFO IN:I OUT:O VDD:B VSS:B
Mm2 OUT IN VSS VSS n_18 W=500.0n L=180n m=1
Mm1 OUT IN VDD VDD p_18 W=1.85u L=180n m=1
.ENDS

************************************************************************
* Library Name: VLSI
* Cell Name:    NAND2
* View Name:    schematic
************************************************************************

.SUBCKT NAND2 A B VDD VOUT VSS
*.PININFO A:I B:I VOUT:O VDD:B VSS:B
MM2 VOUT B VDD VDD p_18 W=1.85u L=180n m=1
MM3 VOUT A VDD VDD p_18 W=1.85u L=180n m=1
MM0 VOUT A net14 VSS n_18 W=1u L=180.00n m=1
MM1 net14 B VSS VSS n_18 W=1u L=180.00n m=1
.ENDS

************************************************************************
* Library Name: VLSI
* Cell Name:    DFFnand
* View Name:    schematic
************************************************************************

.SUBCKT DFFnand CLK D Q QM Qbar A B clkinv VDD VSS
*.PININFO CLK:I D:I Q:O QM:O Qbar:O VDD:B VSS:B
XI9 CLK clkinv VDD VSS / inv
XI8 clkinv net13 VDD VSS / inv
XI7 QM net13 VDD net22 VSS / NAND2
XI6 net22 net13 VDD net23 VSS / NAND2
XI5 net22 Qbar VDD Q VSS / NAND2
XI4 Q net23 VDD Qbar VSS / NAND2
XI3 QM B VDD net41 VSS / NAND2
XI2 A net41 VDD QM VSS / NAND2
XI1 A clkinv VDD B VSS / NAND2
XI0 D clkinv VDD A VSS / NAND2
.ENDS

