* File: RIS.pex.spi
* Created: Fri Dec 27 02:29:37 2024
* Program "Calibre xRC"
* Version "v2016.4_15.11"
* 
.include "RIS.pex.spi.pex"
.subckt RIS  CLK RST VDD VSS M1 M0 CH3 CH2 CH1 CH0
* 
* CH1	CH1
* CH0	CH0
* CH2	CH2
* CH3	CH3
* M1	M1
* CLK	CLK
* M0	M0
* VDD	VDD
* VSS	VSS
* RST	RST
mXI25/XI4/MM2 N_XI25/XI4/NET14_XI25/XI4/MM2_d N_XI25/XI4/NET22_XI25/XI4/MM2_g
+ N_VSS_XI25/XI4/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI4/MM3 N_LFSR10_XI25/XI4/MM3_d N_LFSR10_BAR_XI25/XI4/MM3_g
+ N_VSS_XI25/XI4/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI4/MM10 N_LFSR10_BAR_XI25/XI4/MM10_d N_CLK_XI25/XI4/MM10_g
+ N_XI25/XI4/NET14_XI25/XI4/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI4/XI10/MM3 N_NET089_XI4/XI10/MM3_d N_NET088_XI4/XI10/MM3_g
+ N_VSS_XI4/XI10/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.5e-13 PD=1.48e-06 PS=1.5e-06
mXI4/XI8/MM0 N_XI4/XI8/NET47_XI4/XI8/MM0_d N_NET089_XI4/XI8/MM0_g
+ N_VSS_XI4/XI8/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI0/MM0 N_XI25/XI0/NET6_XI25/XI0/MM0_d N_LFSR10_XI25/XI0/MM0_g
+ N_VSS_XI25/XI0/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI4/MM1 N_XI25/XI4/NET10_XI25/XI4/MM1_d N_CLK_XI25/XI4/MM1_g
+ N_VSS_XI25/XI4/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI4/XI8/MM11 N_XI4/NET031_XI4/XI8/MM11_d N_RSTO_XI4/XI8/MM11_g
+ N_VSS_XI4/XI8/MM11_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=7.5e-07
+ AD=3.675e-13 AS=1.9125e-13 PD=1.73e-06 PS=5.1e-07
mXI18/XI2/XI1/MM0 N_XI18/NET40_XI18/XI2/XI1/MM0_d N_LFSR1_XI18/XI2/XI1/MM0_g
+ N_NET071_XI18/XI2/XI1/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI3/XI1/MM0 N_XI18/NET23_XI18/XI3/XI1/MM0_d N_LFSR1_XI18/XI3/XI1/MM0_g
+ N_NET070_XI18/XI3/XI1/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI4/MM9 N_XI25/XI4/NET22_XI25/XI4/MM9_d N_XI25/XI4/NET6_XI25/XI4/MM9_g
+ N_XI25/XI4/NET10_XI25/XI4/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI4/XI8/MM9 N_XI4/XI8/NET31_XI4/XI8/MM9_d N_XI4/XI8/NET47_XI4/XI8/MM9_g
+ N_XI4/XI8/NET43_XI4/XI8/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI4/XI8/MM11@2 N_XI4/NET031_XI4/XI8/MM11@2_d N_RSTO_XI4/XI8/MM11@2_g
+ N_VSS_XI4/XI8/MM11@2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=7.5e-07
+ AD=3.675e-13 AS=1.9125e-13 PD=1.73e-06 PS=5.1e-07
mXI4/XI8/MM1 N_XI4/XI8/NET43_XI4/XI8/MM1_d N_CLK_XI4/XI8/MM1_g
+ N_VSS_XI4/XI8/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.55e-13 PD=2.5e-07 PS=1.52e-06
mXI25/XI0/MM9 N_XI25/XI0/NET22_XI25/XI0/MM9_d N_XI25/XI0/NET6_XI25/XI0/MM9_g
+ N_XI25/XI0/NET10_XI25/XI0/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI18/XI2/XI2/MM0 N_XI18/NET16_XI18/XI2/XI2/MM0_d N_LFSR1_BAR_XI18/XI2/XI2/MM0_g
+ N_NET071_XI18/XI2/XI2/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI3/XI2/MM0 N_XI18/NET47_XI18/XI3/XI2/MM0_d N_LFSR1_BAR_XI18/XI3/XI2/MM0_g
+ N_NET070_XI18/XI3/XI2/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI0/MM1 N_XI25/XI0/NET10_XI25/XI0/MM1_d N_CLK_XI25/XI0/MM1_g
+ N_VSS_XI25/XI0/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI4/MM0 N_XI25/XI4/NET6_XI25/XI4/MM0_d N_LFSR9_XI25/XI4/MM0_g
+ N_VSS_XI25/XI4/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI4/XI10/MM10 N_NET088_XI4/XI10/MM10_d N_CLK_XI4/XI10/MM10_g
+ N_XI4/XI10/NET16_XI4/XI10/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI4/XI10/MM2 N_XI4/XI10/NET16_XI4/XI10/MM2_d N_XI4/XI10/NET24_XI4/XI10/MM2_g
+ N_VSS_XI4/XI10/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI4/XI8/MM2 N_XI4/XI8/NET39_XI4/XI8/MM2_d N_XI4/XI8/NET31_XI4/XI8/MM2_g
+ N_VSS_XI4/XI8/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI0/MM10 N_LFSR1_BAR_XI25/XI0/MM10_d N_CLK_XI25/XI0/MM10_g
+ N_XI25/XI0/NET14_XI25/XI0/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI4/XI8/MM10 N_XI4/NET031_XI4/XI8/MM10_d N_CLK_XI4/XI8/MM10_g
+ N_XI4/XI8/NET39_XI4/XI8/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.9e-13 AS=6.25e-14 PD=1.66e-06 PS=2.5e-07
mXI25/XI5/MM3 N_LFSR9_XI25/XI5/MM3_d N_LFSR9_BAR_XI25/XI5/MM3_g
+ N_VSS_XI25/XI5/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI0/MM2 N_XI25/XI0/NET14_XI25/XI0/MM2_d N_XI25/XI0/NET22_XI25/XI0/MM2_g
+ N_VSS_XI25/XI0/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI18/XI1/MM3 N_XI18/NET12_XI18/XI1/MM3_d N_XI18/NET16_XI18/XI1/MM3_g
+ N_VSS_XI18/XI1/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI4/MM3 N_XI18/NET19_XI18/XI4/MM3_d N_XI18/NET23_XI18/XI4/MM3_g
+ N_VSS_XI18/XI4/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI4/XI10/MM1 N_XI4/XI10/NET12_XI4/XI10/MM1_d N_CLK_XI4/XI10/MM1_g
+ N_VSS_XI4/XI10/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI4/XI10/MM9 N_XI4/XI10/NET24_XI4/XI10/MM9_d N_XI4/XI10/NET8_XI4/XI10/MM9_g
+ N_XI4/XI10/NET12_XI4/XI10/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI4/XI8/MM3 N_NET087_XI4/XI8/MM3_d N_XI4/NET031_XI4/XI8/MM3_g
+ N_VSS_XI4/XI8/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI5/MM2 N_XI25/XI5/NET14_XI25/XI5/MM2_d N_XI25/XI5/NET22_XI25/XI5/MM2_g
+ N_VSS_XI25/XI5/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI0/MM3 N_LFSR1_XI25/XI0/MM3_d N_LFSR1_BAR_XI25/XI0/MM3_g
+ N_VSS_XI25/XI0/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI5/MM10 N_LFSR9_BAR_XI25/XI5/MM10_d N_CLK_XI25/XI5/MM10_g
+ N_XI25/XI5/NET14_XI25/XI5/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI4/XI10/MM0 N_XI4/XI10/NET8_XI4/XI10/MM0_d N_XI4/NET031_XI4/XI10/MM0_g
+ N_VSS_XI4/XI10/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI1/MM10 N_XI18/NET16_XI18/XI1/MM10_d N_CLK_XI18/XI1/MM10_g
+ N_XI18/XI1/NET16_XI18/XI1/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI18/XI4/MM10 N_XI18/NET23_XI18/XI4/MM10_d N_CLK_XI18/XI4/MM10_g
+ N_XI18/XI4/NET16_XI18/XI4/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI25/XI5/MM1 N_XI25/XI5/NET10_XI25/XI5/MM1_d N_CLK_XI25/XI5/MM1_g
+ N_VSS_XI25/XI5/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI6/MM0 N_XI25/XI6/NET47_XI25/XI6/MM0_d N_LFSR1_XI25/XI6/MM0_g
+ N_VSS_XI25/XI6/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI1/MM2 N_XI18/XI1/NET16_XI18/XI1/MM2_d N_XI18/XI1/NET24_XI18/XI1/MM2_g
+ N_VSS_XI18/XI1/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI18/XI4/MM2 N_XI18/XI4/NET16_XI18/XI4/MM2_d N_XI18/XI4/NET24_XI18/XI4/MM2_g
+ N_VSS_XI18/XI4/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI23/MM0 N_RST_XI23/MM0_d N_CLK_XI23/MM0_g N_RSTO_XI23/MM0_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI25/XI5/MM9 N_XI25/XI5/NET22_XI25/XI5/MM9_d N_XI25/XI5/NET6_XI25/XI5/MM9_g
+ N_XI25/XI5/NET10_XI25/XI5/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI18/XI1/MM1 N_XI18/XI1/NET12_XI18/XI1/MM1_d N_CLK_XI18/XI1/MM1_g
+ N_VSS_XI18/XI1/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI18/XI4/MM1 N_XI18/XI4/NET12_XI18/XI4/MM1_d N_CLK_XI18/XI4/MM1_g
+ N_VSS_XI18/XI4/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI5/MM0 N_XI25/XI5/NET6_XI25/XI5/MM0_d N_LFSR8_XI25/XI5/MM0_g
+ N_VSS_XI25/XI5/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI6/MM9 N_XI25/XI6/NET31_XI25/XI6/MM9_d N_XI25/XI6/NET47_XI25/XI6/MM9_g
+ N_XI25/XI6/NET43_XI25/XI6/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI24/Mm2 N_CLKBAR_XI24/Mm2_d N_CLK_XI24/Mm2_g N_VSS_XI24/Mm2_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=2.5e-07 AD=2.509e-13 AS=2.509e-13
+ PD=1.87e-06 PS=1.87e-06
mXI18/XI1/MM9 N_XI18/XI1/NET24_XI18/XI1/MM9_d N_XI18/XI1/NET8_XI18/XI1/MM9_g
+ N_XI18/XI1/NET12_XI18/XI1/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI18/XI4/MM9 N_XI18/XI4/NET24_XI18/XI4/MM9_d N_XI18/XI4/NET8_XI18/XI4/MM9_g
+ N_XI18/XI4/NET12_XI18/XI4/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI25/XI6/MM1 N_XI25/XI6/NET43_XI25/XI6/MM1_d N_CLK_XI25/XI6/MM1_g
+ N_VSS_XI25/XI6/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=3.525e-13 PD=2.5e-07 PS=1.91e-06
mXI13/Mm2 N_RSTOBAR_XI13/Mm2_d N_RSTO_XI13/Mm2_g N_VSS_XI13/Mm2_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=2.5e-07 AD=2.509e-13 AS=2.509e-13
+ PD=1.87e-06 PS=1.87e-06
mXI25/XI1/MM3 N_LFSR8_XI25/XI1/MM3_d N_LFSR8_BAR_XI25/XI1/MM3_g
+ N_VSS_XI25/XI1/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI1/MM0 N_XI18/XI1/NET8_XI18/XI1/MM0_d N_XI18/PREBIT0_XI18/XI1/MM0_g
+ N_VSS_XI18/XI1/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI4/MM0 N_XI18/XI4/NET8_XI18/XI4/MM0_d N_XI18/PREBIT1_XI18/XI4/MM0_g
+ N_VSS_XI18/XI4/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI6/MM2 N_XI25/XI6/NET39_XI25/XI6/MM2_d N_XI25/XI6/NET31_XI25/XI6/MM2_g
+ N_VSS_XI25/XI6/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI6/MM10 N_LFSR2_BAR_XI25/XI6/MM10_d N_CLK_XI25/XI6/MM10_g
+ N_XI25/XI6/NET39_XI25/XI6/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.9e-13 AS=6.25e-14 PD=1.66e-06 PS=2.5e-07
mXI25/XI1/MM2 N_XI25/XI1/NET14_XI25/XI1/MM2_d N_XI25/XI1/NET22_XI25/XI1/MM2_g
+ N_VSS_XI25/XI1/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI17/XI7/MM3 N_XI17/A0_XI17/XI7/MM3_d N_XI17/A0BAR_XI17/XI7/MM3_g
+ N_VSS_XI17/XI7/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI6/MM3 N_XI17/A1_XI17/XI6/MM3_d N_XI17/A1BAR_XI17/XI6/MM3_g
+ N_VSS_XI17/XI6/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI1/MM10 N_LFSR8_BAR_XI25/XI1/MM10_d N_CLK_XI25/XI1/MM10_g
+ N_XI25/XI1/NET14_XI25/XI1/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI18/XI6/MM11 N_XI18/NET40_XI18/XI6/MM11_d N_RSTO_XI18/XI6/MM11_g
+ N_VSS_XI18/XI6/MM11_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI18/XI9/MM11 N_XI18/NET47_XI18/XI9/MM11_d N_RSTO_XI18/XI9/MM11_g
+ N_VSS_XI18/XI9/MM11_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI25/XI6/MM3 N_LFSR2_XI25/XI6/MM3_d N_LFSR2_BAR_XI25/XI6/MM3_g
+ N_VSS_XI25/XI6/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI1/MM1 N_XI25/XI1/NET10_XI25/XI1/MM1_d N_CLK_XI25/XI1/MM1_g
+ N_VSS_XI25/XI1/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI1/MM9 N_XI25/XI1/NET22_XI25/XI1/MM9_d N_XI25/XI1/NET6_XI25/XI1/MM9_g
+ N_XI25/XI1/NET10_XI25/XI1/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI18/XI6/MM3 N_XI18/PREBIT0_XI18/XI6/MM3_d N_XI18/NET40_XI18/XI6/MM3_g
+ N_VSS_XI18/XI6/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI9/MM3 N_XI18/PREBIT1_XI18/XI9/MM3_d N_XI18/NET47_XI18/XI9/MM3_g
+ N_VSS_XI18/XI9/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI7/MM10 N_XI17/A0BAR_XI17/XI7/MM10_d N_CLK_XI17/XI7/MM10_g
+ N_XI17/XI7/NET16_XI17/XI7/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI17/XI6/MM10 N_XI17/A1BAR_XI17/XI6/MM10_d N_CLK_XI17/XI6/MM10_g
+ N_XI17/XI6/NET16_XI17/XI6/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI25/XI6/MM11 N_LFSR2_BAR_XI25/XI6/MM11_d N_RST_XI25/XI6/MM11_g
+ N_VSS_XI25/XI6/MM11_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=1.5e-06
+ AD=7.35e-13 AS=7.35e-13 PD=2.48e-06 PS=2.48e-06
mXI17/XI7/MM2 N_XI17/XI7/NET16_XI17/XI7/MM2_d N_XI17/XI7/NET24_XI17/XI7/MM2_g
+ N_VSS_XI17/XI7/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI17/XI6/MM2 N_XI17/XI6/NET16_XI17/XI6/MM2_d N_XI17/XI6/NET24_XI17/XI6/MM2_g
+ N_VSS_XI17/XI6/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI1/MM0 N_XI25/XI1/NET6_XI25/XI1/MM0_d N_LFSR7_XI25/XI1/MM0_g
+ N_VSS_XI25/XI1/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI6/MM10 N_XI18/NET40_XI18/XI6/MM10_d N_CLK_XI18/XI6/MM10_g
+ N_XI18/XI6/NET39_XI18/XI6/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.9e-13 AS=6.25e-14 PD=1.66e-06 PS=2.5e-07
mXI18/XI9/MM10 N_XI18/NET47_XI18/XI9/MM10_d N_CLK_XI18/XI9/MM10_g
+ N_XI18/XI9/NET39_XI18/XI9/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.9e-13 AS=6.25e-14 PD=1.66e-06 PS=2.5e-07
mXI18/XI6/MM2 N_XI18/XI6/NET39_XI18/XI6/MM2_d N_XI18/XI6/NET31_XI18/XI6/MM2_g
+ N_VSS_XI18/XI6/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI18/XI9/MM2 N_XI18/XI9/NET39_XI18/XI9/MM2_d N_XI18/XI9/NET31_XI18/XI9/MM2_g
+ N_VSS_XI18/XI9/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI3/MM3 N_LFSR7_XI25/XI3/MM3_d N_LFSR7_BAR_XI25/XI3/MM3_g
+ N_VSS_XI25/XI3/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI7/MM1 N_XI17/XI7/NET12_XI17/XI7/MM1_d N_CLK_XI17/XI7/MM1_g
+ N_VSS_XI17/XI7/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI17/XI6/MM1 N_XI17/XI6/NET12_XI17/XI6/MM1_d N_CLK_XI17/XI6/MM1_g
+ N_VSS_XI17/XI6/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI18/MM0 N_XI25/XI18/NET6_XI25/XI18/MM0_d N_LFSR2_XI25/XI18/MM0_g
+ N_VSS_XI25/XI18/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI7/MM9 N_XI17/XI7/NET24_XI17/XI7/MM9_d N_XI17/XI7/NET8_XI17/XI7/MM9_g
+ N_XI17/XI7/NET12_XI17/XI7/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI17/XI6/MM9 N_XI17/XI6/NET24_XI17/XI6/MM9_d N_XI17/XI6/NET8_XI17/XI6/MM9_g
+ N_XI17/XI6/NET12_XI17/XI6/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI25/XI3/MM2 N_XI25/XI3/NET14_XI25/XI3/MM2_d N_XI25/XI3/NET22_XI25/XI3/MM2_g
+ N_VSS_XI25/XI3/MM2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI18/XI6/MM1 N_XI18/XI6/NET43_XI18/XI6/MM1_d N_CLK_XI18/XI6/MM1_g
+ N_VSS_XI18/XI6/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=3.525e-13 PD=2.5e-07 PS=1.91e-06
mXI18/XI9/MM1 N_XI18/XI9/NET43_XI18/XI9/MM1_d N_CLK_XI18/XI9/MM1_g
+ N_VSS_XI18/XI9/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=3.525e-13 PD=2.5e-07 PS=1.91e-06
mXI25/XI18/MM9 N_XI25/XI18/NET22_XI25/XI18/MM9_d
+ N_XI25/XI18/NET6_XI25/XI18/MM9_g N_XI25/XI18/NET10_XI25/XI18/MM9_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=6.25e-14
+ PD=1.48e-06 PS=2.5e-07
mXI25/XI3/MM10 N_LFSR7_BAR_XI25/XI3/MM10_d N_CLK_XI25/XI3/MM10_g
+ N_XI25/XI3/NET14_XI25/XI3/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI17/XI7/MM0 N_XI17/XI7/NET8_XI17/XI7/MM0_d N_NET083_XI17/XI7/MM0_g
+ N_VSS_XI17/XI7/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI6/MM0 N_XI17/XI6/NET8_XI17/XI6/MM0_d N_NET082_XI17/XI6/MM0_g
+ N_VSS_XI17/XI6/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI6/MM9 N_XI18/XI6/NET31_XI18/XI6/MM9_d N_XI18/XI6/NET47_XI18/XI6/MM9_g
+ N_XI18/XI6/NET43_XI18/XI6/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI18/XI9/MM9 N_XI18/XI9/NET31_XI18/XI9/MM9_d N_XI18/XI9/NET47_XI18/XI9/MM9_g
+ N_XI18/XI9/NET43_XI18/XI9/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI25/XI18/MM1 N_XI25/XI18/NET10_XI25/XI18/MM1_d N_CLK_XI25/XI18/MM1_g
+ N_VSS_XI25/XI18/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI3/MM1 N_XI25/XI3/NET10_XI25/XI3/MM1_d N_CLK_XI25/XI3/MM1_g
+ N_VSS_XI25/XI3/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI18/MM10 N_LFSR3_BAR_XI25/XI18/MM10_d N_CLK_XI25/XI18/MM10_g
+ N_XI25/XI18/NET14_XI25/XI18/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI17/XI1/XI2/MM0 N_XI17/NET13_XI17/XI1/XI2/MM0_d N_LFSR7_BAR_XI17/XI1/XI2/MM0_g
+ N_NET082_XI17/XI1/XI2/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI4/XI2/MM0 N_XI17/NET024_XI17/XI4/XI2/MM0_d N_LFSR7_XI17/XI4/XI2/MM0_g
+ N_NET083_XI17/XI4/XI2/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI3/MM9 N_XI25/XI3/NET22_XI25/XI3/MM9_d N_XI25/XI3/NET6_XI25/XI3/MM9_g
+ N_XI25/XI3/NET10_XI25/XI3/MM9_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI18/XI6/MM0 N_XI18/XI6/NET47_XI18/XI6/MM0_d N_NET071_XI18/XI6/MM0_g
+ N_VSS_XI18/XI6/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI9/MM0 N_XI18/XI9/NET47_XI18/XI9/MM0_d N_NET070_XI18/XI9/MM0_g
+ N_VSS_XI18/XI9/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI18/MM2 N_XI25/XI18/NET14_XI25/XI18/MM2_d
+ N_XI25/XI18/NET22_XI25/XI18/MM2_g N_VSS_XI25/XI18/MM2_s N_VSS_XI25/XI4/MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=6.25e-14 AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI17/XI1/XI1/MM0 N_XI17/A1BAR_XI17/XI1/XI1/MM0_d N_LFSR7_XI17/XI1/XI1/MM0_g
+ N_NET082_XI17/XI1/XI1/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI4/XI1/MM0 N_XI17/A0BAR_XI17/XI4/XI1/MM0_d N_LFSR7_BAR_XI17/XI4/XI1/MM0_g
+ N_NET083_XI17/XI4/XI1/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI3/MM0 N_XI25/XI3/NET6_XI25/XI3/MM0_d N_LFSR6_XI25/XI3/MM0_g
+ N_VSS_XI25/XI3/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI18/MM3 N_LFSR3_XI25/XI18/MM3_d N_LFSR3_BAR_XI25/XI18/MM3_g
+ N_VSS_XI25/XI18/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI0/XI2/MM0 N_NET071_XI5/XI0/XI0/XI2/MM0_d
+ N_M0_BAR_XI5/XI0/XI0/XI2/MM0_g N_XI5/XI0/NET40_XI5/XI0/XI0/XI2/MM0_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI0/XI1/MM0 N_NET089_XI5/XI0/XI0/XI1/MM0_d N_M0_XI5/XI0/XI0/XI1/MM0_g
+ N_XI5/XI0/NET40_XI5/XI0/XI0/XI1/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI7/XI1/MM0 N_NET087_XI5/XI0/XI7/XI1/MM0_d N_M0_XI5/XI0/XI7/XI1/MM0_g
+ N_XI5/XI0/NET33_XI5/XI0/XI7/XI1/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI7/XI2/MM0 N_NET070_XI5/XI0/XI7/XI2/MM0_d
+ N_M0_BAR_XI5/XI0/XI7/XI2/MM0_g N_XI5/XI0/NET33_XI5/XI0/XI7/XI2/MM0_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI25/XI14/MM3 N_LFSR6_XI25/XI14/MM3_d N_LFSR6_BAR_XI25/XI14/MM3_g
+ N_VSS_XI25/XI14/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI2/XI2/MM0 N_LFSR3_BAR_XI25/XI2/XI2/MM0_d N_LFSR10_XI25/XI2/XI2/MM0_g
+ N_XI25/NET62_XI25/XI2/XI2/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI2/XI2/MM0 N_XI17/A1_XI17/XI2/XI2/MM0_d N_LFSR5_BAR_XI17/XI2/XI2/MM0_g
+ N_XI17/NET13_XI17/XI2/XI2/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI3/XI2/MM0 N_XI17/A0_XI17/XI3/XI2/MM0_d N_LFSR5_BAR_XI17/XI3/XI2/MM0_g
+ N_XI17/NET024_XI17/XI3/XI2/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI14/MM2 N_XI25/XI14/NET14_XI25/XI14/MM2_d
+ N_XI25/XI14/NET22_XI25/XI14/MM2_g N_VSS_XI25/XI14/MM2_s N_VSS_XI25/XI4/MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=6.25e-14 AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI2/XI3/MM0 N_LFSR3_XI25/XI2/XI3/MM0_d N_LFSR10_BAR_XI25/XI2/XI3/MM0_g
+ N_XI25/NET62_XI25/XI2/XI3/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI14/MM10 N_LFSR6_BAR_XI25/XI14/MM10_d N_CLK_XI25/XI14/MM10_g
+ N_XI25/XI14/NET14_XI25/XI14/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI17/XI2/XI1/MM0 N_LFSR6_XI17/XI2/XI1/MM0_d N_LFSR5_XI17/XI2/XI1/MM0_g
+ N_XI17/NET13_XI17/XI2/XI1/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI3/XI1/MM0 N_LFSR6_XI17/XI3/XI1/MM0_d N_LFSR5_XI17/XI3/XI1/MM0_g
+ N_XI17/NET024_XI17/XI3/XI1/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI16/MM0 N_XI25/XI16/NET6_XI25/XI16/MM0_d N_XI25/NET62_XI25/XI16/MM0_g
+ N_VSS_XI25/XI16/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI14/MM1 N_XI25/XI14/NET10_XI25/XI14/MM1_d N_CLK_XI25/XI14/MM1_g
+ N_VSS_XI25/XI14/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI14/MM9 N_XI25/XI14/NET22_XI25/XI14/MM9_d
+ N_XI25/XI14/NET6_XI25/XI14/MM9_g N_XI25/XI14/NET10_XI25/XI14/MM9_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=6.25e-14
+ PD=1.48e-06 PS=2.5e-07
mXI5/XI0/XI2/XI2/MM0 N_XI5/XI0/NET54_XI5/XI0/XI2/XI2/MM0_d
+ N_M1_BAR_XI5/XI0/XI2/XI2/MM0_g N_XI5/NET64_XI5/XI0/XI2/XI2/MM0_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI2/XI1/MM0 N_XI5/XI0/NET40_XI5/XI0/XI2/XI1/MM0_d
+ N_M1_XI5/XI0/XI2/XI1/MM0_g N_XI5/NET64_XI5/XI0/XI2/XI1/MM0_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI8/XI1/MM0 N_XI5/XI0/NET33_XI5/XI0/XI8/XI1/MM0_d
+ N_M1_XI5/XI0/XI8/XI1/MM0_g N_XI5/NET63_XI5/XI0/XI8/XI1/MM0_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI8/XI2/MM0 N_XI5/XI0/NET19_XI5/XI0/XI8/XI2/MM0_d
+ N_M1_BAR_XI5/XI0/XI8/XI2/MM0_g N_XI5/NET63_XI5/XI0/XI8/XI2/MM0_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI25/XI16/MM9 N_XI25/XI16/NET22_XI25/XI16/MM9_d
+ N_XI25/XI16/NET6_XI25/XI16/MM9_g N_XI25/XI16/NET10_XI25/XI16/MM9_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=6.25e-14
+ PD=1.48e-06 PS=2.5e-07
mXI25/XI16/MM1 N_XI25/XI16/NET10_XI25/XI16/MM1_d N_CLK_XI25/XI16/MM1_g
+ N_VSS_XI25/XI16/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI5/XI0/XI9/XI2/MM0 N_LFSR8_XI5/XI0/XI9/XI2/MM0_d
+ N_M0_BAR_XI5/XI0/XI9/XI2/MM0_g N_XI5/XI0/NET19_XI5/XI0/XI9/XI2/MM0_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI9/XI1/MM0 N_NET082_XI5/XI0/XI9/XI1/MM0_d N_M0_XI5/XI0/XI9/XI1/MM0_g
+ N_XI5/XI0/NET19_XI5/XI0/XI9/XI1/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI1/XI1/MM0 N_NET083_XI5/XI0/XI1/XI1/MM0_d N_M0_XI5/XI0/XI1/XI1/MM0_g
+ N_XI5/XI0/NET54_XI5/XI0/XI1/XI1/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI1/XI2/MM0 N_LFSR3_XI5/XI0/XI1/XI2/MM0_d
+ N_M0_BAR_XI5/XI0/XI1/XI2/MM0_g N_XI5/XI0/NET54_XI5/XI0/XI1/XI2/MM0_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI25/XI14/MM0 N_XI25/XI14/NET6_XI25/XI14/MM0_d N_LFSR5_XI25/XI14/MM0_g
+ N_VSS_XI25/XI14/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI16/MM10 N_LFSR4_BAR_XI25/XI16/MM10_d N_CLK_XI25/XI16/MM10_g
+ N_XI25/XI16/NET14_XI25/XI16/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI25/XI15/MM3 N_LFSR5_XI25/XI15/MM3_d N_LFSR5_BAR_XI25/XI15/MM3_g
+ N_VSS_XI25/XI15/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI16/MM2 N_XI25/XI16/NET14_XI25/XI16/MM2_d
+ N_XI25/XI16/NET22_XI25/XI16/MM2_g N_VSS_XI25/XI16/MM2_s N_VSS_XI25/XI4/MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=6.25e-14 AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI15/MM2 N_XI25/XI15/NET14_XI25/XI15/MM2_d
+ N_XI25/XI15/NET22_XI25/XI15/MM2_g N_VSS_XI25/XI15/MM2_s N_VSS_XI25/XI4/MM2_b
+ N_18 L=1.8e-07 W=5e-07 AD=6.25e-14 AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI16/MM3 N_LFSR4_XI25/XI16/MM3_d N_LFSR4_BAR_XI25/XI16/MM3_g
+ N_VSS_XI25/XI16/MM3_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI15/MM10 N_LFSR5_BAR_XI25/XI15/MM10_d N_CLK_XI25/XI15/MM10_g
+ N_XI25/XI15/NET14_XI25/XI15/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=6.25e-14 PD=1.48e-06 PS=2.5e-07
mXI5/XI2/Mm2 N_XI5/NET42_XI5/XI2/Mm2_d N_XI5/NET64_XI5/XI2/Mm2_g
+ N_VSS_XI5/XI2/Mm2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=2.5e-07 AD=2.509e-13
+ AS=2.509e-13 PD=1.87e-06 PS=1.87e-06
mXI5/XI3/Mm2 N_XI5/NET38_XI5/XI3/Mm2_d N_XI5/NET63_XI5/XI3/Mm2_g
+ N_VSS_XI5/XI3/Mm2_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=2.5e-07 AD=2.509e-13
+ AS=2.509e-13 PD=1.87e-06 PS=1.87e-06
mXI7/Mm2 N_M0_BAR_XI7/Mm2_d N_M0_XI7/Mm2_g N_VSS_XI7/Mm2_s N_VSS_XI25/XI4/MM2_b
+ N_18 L=1.8e-07 W=2.5e-07 AD=2.509e-13 AS=2.509e-13 PD=1.87e-06 PS=1.87e-06
mXI8/Mm2 N_M1_BAR_XI8/Mm2_d N_M1_XI8/Mm2_g N_VSS_XI8/Mm2_s N_VSS_XI25/XI4/MM2_b
+ N_18 L=1.8e-07 W=2.5e-07 AD=2.509e-13 AS=2.509e-13 PD=1.87e-06 PS=1.87e-06
mXI25/XI15/MM1 N_XI25/XI15/NET10_XI25/XI15/MM1_d N_CLK_XI25/XI15/MM1_g
+ N_VSS_XI25/XI15/MM1_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=6.25e-14
+ AS=2.45e-13 PD=2.5e-07 PS=1.48e-06
mXI25/XI15/MM9 N_XI25/XI15/NET22_XI25/XI15/MM9_d
+ N_XI25/XI15/NET6_XI25/XI15/MM9_g N_XI25/XI15/NET10_XI25/XI15/MM9_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=6.25e-14
+ PD=1.48e-06 PS=2.5e-07
mXI5/XI1/MM15 N_VSS_XI5/XI1/MM15_d N_XI5/NET42_XI5/XI1/MM15_g
+ N_CH3_XI5/XI1/MM15_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=2.5e-07
+ AD=2.509e-13 AS=1.4045e-13 PD=1.87e-06 PS=9.3e-07
mXI5/XI1/MM0 N_VSS_XI5/XI1/MM0_d N_XI5/NET64_XI5/XI1/MM0_g N_CH0_XI5/XI1/MM0_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=2.5e-07 AD=2.509e-13 AS=1.4045e-13
+ PD=1.87e-06 PS=9.3e-07
mXI5/XI1/MM7 N_VSS_XI5/XI1/MM7_d N_XI5/NET42_XI5/XI1/MM7_g N_CH1_XI5/XI1/MM7_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=2.5e-07 AD=2.509e-13 AS=1.4045e-13
+ PD=1.87e-06 PS=9.3e-07
mXI5/XI1/MM10 N_VSS_XI5/XI1/MM10_d N_XI5/NET64_XI5/XI1/MM10_g
+ N_CH2_XI5/XI1/MM10_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=2.5e-07
+ AD=2.509e-13 AS=1.4045e-13 PD=1.87e-06 PS=9.3e-07
mXI5/XI1/MM14 N_VSS_XI5/XI1/MM14_d N_XI5/NET38_XI5/XI1/MM14_g
+ N_CH3_XI5/XI1/MM14_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=2.5e-07
+ AD=2.509e-13 AS=1.4045e-13 PD=1.87e-06 PS=9.3e-07
mXI5/XI1/MM1 N_VSS_XI5/XI1/MM1_d N_XI5/NET63_XI5/XI1/MM1_g N_CH0_XI5/XI1/MM1_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=2.5e-07 AD=2.509e-13 AS=1.4045e-13
+ PD=1.87e-06 PS=9.3e-07
mXI5/XI1/MM6 N_VSS_XI5/XI1/MM6_d N_XI5/NET63_XI5/XI1/MM6_g N_CH1_XI5/XI1/MM6_s
+ N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=2.5e-07 AD=2.509e-13 AS=1.4045e-13
+ PD=1.87e-06 PS=9.3e-07
mXI5/XI1/MM11 N_VSS_XI5/XI1/MM11_d N_XI5/NET38_XI5/XI1/MM11_g
+ N_CH2_XI5/XI1/MM11_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=2.5e-07
+ AD=2.509e-13 AS=1.4045e-13 PD=1.87e-06 PS=9.3e-07
mXI25/XI15/MM0 N_XI25/XI15/NET6_XI25/XI15/MM0_d N_LFSR4_XI25/XI15/MM0_g
+ N_VSS_XI25/XI15/MM0_s N_VSS_XI25/XI4/MM2_b N_18 L=1.8e-07 W=5e-07 AD=2.45e-13
+ AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI4/MM7 N_LFSR10_BAR_XI25/XI4/MM7_d N_XI25/XI4/NET22_XI25/XI4/MM7_g
+ N_VDD_XI25/XI4/MM7_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI4/MM8 N_LFSR10_XI25/XI4/MM8_d N_LFSR10_BAR_XI25/XI4/MM8_g
+ N_VDD_XI25/XI4/MM8_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI4/XI10/MM8 N_NET089_XI4/XI10/MM8_d N_NET088_XI4/XI10/MM8_g
+ N_VDD_XI4/XI10/MM8_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI4/XI8/MM5 N_XI4/XI8/NET26_XI4/XI8/MM5_d N_NET089_XI4/XI8/MM5_g
+ N_VDD_XI4/XI8/MM5_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=7e-07 AD=8.75e-14
+ AS=3.43e-13 PD=2.5e-07 PS=1.68e-06
mXI4/XI8/MM4 N_XI4/XI8/NET47_XI4/XI8/MM4_d N_CLK_XI4/XI8/MM4_g
+ N_XI4/XI8/NET26_XI4/XI8/MM4_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=7e-07
+ AD=4.095e-13 AS=8.75e-14 PD=1.87e-06 PS=2.5e-07
mXI25/XI0/MM5 N_XI25/XI0/NET33_XI25/XI0/MM5_d N_LFSR10_XI25/XI0/MM5_g
+ N_VDD_XI25/XI0/MM5_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06 AD=2.25e-13
+ AS=8.82e-13 PD=2.5e-07 PS=2.78e-06
mXI25/XI4/MM6 N_XI25/XI4/NET22_XI25/XI4/MM6_d N_CLK_XI25/XI4/MM6_g
+ N_VDD_XI25/XI4/MM6_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI0/MM4 N_XI25/XI0/NET6_XI25/XI0/MM4_d N_CLK_XI25/XI0/MM4_g
+ N_XI25/XI0/NET33_XI25/XI0/MM4_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=2.25e-13 PD=2.78e-06 PS=2.5e-07
mXI4/XI10/MM11 N_NET088_XI4/XI10/MM11_d N_RSTOBAR_XI4/XI10/MM11_g
+ N_VDD_XI4/XI10/MM11_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI18/XI2/XI1/MM1 N_XI18/NET40_XI18/XI2/XI1/MM1_d N_LFSR1_BAR_XI18/XI2/XI1/MM1_g
+ N_NET071_XI18/XI2/XI1/MM1_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI3/XI1/MM1 N_XI18/NET23_XI18/XI3/XI1/MM1_d N_LFSR1_BAR_XI18/XI3/XI1/MM1_g
+ N_NET070_XI18/XI3/XI1/MM1_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI4/XI8/MM6 N_XI4/XI8/NET31_XI4/XI8/MM6_d N_CLK_XI4/XI8/MM6_g
+ N_VDD_XI4/XI8/MM6_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=4.935e-13 PD=1.68e-06 PS=2.11e-06
mXI18/XI2/XI2/MM1 N_XI18/NET16_XI18/XI2/XI2/MM1_d N_LFSR1_XI18/XI2/XI2/MM1_g
+ N_NET071_XI18/XI2/XI2/MM1_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI18/XI3/XI2/MM1 N_XI18/NET47_XI18/XI3/XI2/MM1_d N_LFSR1_XI18/XI3/XI2/MM1_g
+ N_NET070_XI18/XI3/XI2/MM1_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI4/MM4 N_XI25/XI4/NET6_XI25/XI4/MM4_d N_CLK_XI25/XI4/MM4_g
+ N_XI25/XI4/NET33_XI25/XI4/MM4_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=2.25e-13 PD=2.78e-06 PS=2.5e-07
mXI25/XI0/MM6 N_XI25/XI0/NET22_XI25/XI0/MM6_d N_CLK_XI25/XI0/MM6_g
+ N_VDD_XI25/XI0/MM6_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI4/MM5 N_XI25/XI4/NET33_XI25/XI4/MM5_d N_LFSR9_XI25/XI4/MM5_g
+ N_VDD_XI25/XI4/MM5_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=2.25e-13
+ AS=8.82e-13 PD=2.5e-07 PS=2.78e-06
mXI4/XI10/MM7 N_NET088_XI4/XI10/MM7_d N_XI4/XI10/NET24_XI4/XI10/MM7_g
+ N_VDD_XI4/XI10/MM7_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.57e-13
+ AS=3.43e-13 PD=1.72e-06 PS=1.68e-06
mXI4/XI8/MM7 N_XI4/NET031_XI4/XI8/MM7_d N_XI4/XI8/NET31_XI4/XI8/MM7_g
+ N_VDD_XI4/XI8/MM7_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=7e-07 AD=7.07e-13
+ AS=3.43e-13 PD=2.72e-06 PS=1.68e-06
mXI25/XI5/MM8 N_LFSR9_XI25/XI5/MM8_d N_LFSR9_BAR_XI25/XI5/MM8_g
+ N_VDD_XI25/XI5/MM8_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI0/MM7 N_LFSR1_BAR_XI25/XI0/MM7_d N_XI25/XI0/NET22_XI25/XI0/MM7_g
+ N_VDD_XI25/XI0/MM7_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI18/XI1/MM8 N_XI18/NET12_XI18/XI1/MM8_d N_XI18/NET16_XI18/XI1/MM8_g
+ N_VDD_XI18/XI1/MM8_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI18/XI4/MM8 N_XI18/NET19_XI18/XI4/MM8_d N_XI18/NET23_XI18/XI4/MM8_g
+ N_VDD_XI18/XI4/MM8_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07 W=7e-07
+ AD=3.43e-13 AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI4/XI10/MM6 N_XI4/XI10/NET24_XI4/XI10/MM6_d N_CLK_XI4/XI10/MM6_g
+ N_VDD_XI4/XI10/MM6_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI4/XI8/MM8 N_NET087_XI4/XI8/MM8_d N_XI4/NET031_XI4/XI8/MM8_g
+ N_VDD_XI4/XI8/MM8_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI25/XI5/MM7 N_LFSR9_BAR_XI25/XI5/MM7_d N_XI25/XI5/NET22_XI25/XI5/MM7_g
+ N_VDD_XI25/XI5/MM7_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI0/MM8 N_LFSR1_XI25/XI0/MM8_d N_LFSR1_BAR_XI25/XI0/MM8_g
+ N_VDD_XI25/XI0/MM8_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI18/XI1/MM11 N_XI18/NET16_XI18/XI1/MM11_d N_RSTOBAR_XI18/XI1/MM11_g
+ N_VDD_XI18/XI1/MM11_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI18/XI4/MM11 N_XI18/NET23_XI18/XI4/MM11_d N_RSTOBAR_XI18/XI4/MM11_g
+ N_VDD_XI18/XI4/MM11_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07 W=7e-07
+ AD=3.43e-13 AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI4/XI10/MM4 N_XI4/XI10/NET8_XI4/XI10/MM4_d N_CLK_XI4/XI10/MM4_g
+ N_XI4/XI10/NET39_XI4/XI10/MM4_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07
+ AD=3.43e-13 AS=8.75e-14 PD=1.68e-06 PS=2.5e-07
mXI4/XI10/MM5 N_XI4/XI10/NET39_XI4/XI10/MM5_d N_XI4/NET031_XI4/XI10/MM5_g
+ N_VDD_XI4/XI10/MM5_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=8.75e-14
+ AS=3.43e-13 PD=2.5e-07 PS=1.68e-06
mXI25/XI5/MM6 N_XI25/XI5/NET22_XI25/XI5/MM6_d N_CLK_XI25/XI5/MM6_g
+ N_VDD_XI25/XI5/MM6_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI6/MM5 N_XI25/XI6/NET26_XI25/XI6/MM5_d N_LFSR1_XI25/XI6/MM5_g
+ N_VDD_XI25/XI6/MM5_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=7e-07 AD=8.75e-14
+ AS=3.43e-13 PD=2.5e-07 PS=1.68e-06
mXI18/XI1/MM7 N_XI18/NET16_XI18/XI1/MM7_d N_XI18/XI1/NET24_XI18/XI1/MM7_g
+ N_VDD_XI18/XI1/MM7_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=6.44e-13
+ AS=3.43e-13 PD=2.54e-06 PS=1.68e-06
mXI18/XI4/MM7 N_XI18/NET23_XI18/XI4/MM7_d N_XI18/XI4/NET24_XI18/XI4/MM7_g
+ N_VDD_XI18/XI4/MM7_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07 W=7e-07
+ AD=6.44e-13 AS=3.43e-13 PD=2.54e-06 PS=1.68e-06
mXI23/MM1 N_RST_XI23/MM1_d N_CLKBAR_XI23/MM1_g N_RSTO_XI23/MM1_s
+ N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06
+ PS=1.48e-06
mXI25/XI6/MM4 N_XI25/XI6/NET47_XI25/XI6/MM4_d N_CLK_XI25/XI6/MM4_g
+ N_XI25/XI6/NET26_XI25/XI6/MM4_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=7e-07
+ AD=4.095e-13 AS=8.75e-14 PD=1.87e-06 PS=2.5e-07
mXI25/XI5/MM4 N_XI25/XI5/NET6_XI25/XI5/MM4_d N_CLK_XI25/XI5/MM4_g
+ N_XI25/XI5/NET33_XI25/XI5/MM4_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=2.25e-13 PD=2.78e-06 PS=2.5e-07
mXI18/XI1/MM6 N_XI18/XI1/NET24_XI18/XI1/MM6_d N_CLK_XI18/XI1/MM6_g
+ N_VDD_XI18/XI1/MM6_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI18/XI4/MM6 N_XI18/XI4/NET24_XI18/XI4/MM6_d N_CLK_XI18/XI4/MM6_g
+ N_VDD_XI18/XI4/MM6_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07 W=7e-07
+ AD=3.43e-13 AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI25/XI5/MM5 N_XI25/XI5/NET33_XI25/XI5/MM5_d N_LFSR8_XI25/XI5/MM5_g
+ N_VDD_XI25/XI5/MM5_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=2.25e-13
+ AS=8.82e-13 PD=2.5e-07 PS=2.78e-06
mXI24/Mm1 N_CLKBAR_XI24/Mm1_d N_CLK_XI24/Mm1_g N_VDD_XI24/Mm1_s
+ N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=3.5e-07 AD=2.629e-13 AS=2.629e-13
+ PD=1.77e-06 PS=1.77e-06
mXI25/XI6/MM6 N_XI25/XI6/NET31_XI25/XI6/MM6_d N_CLK_XI25/XI6/MM6_g
+ N_VDD_XI25/XI6/MM6_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=4.935e-13 PD=1.68e-06 PS=2.11e-06
mXI13/Mm1 N_RSTOBAR_XI13/Mm1_d N_RSTO_XI13/Mm1_g N_VDD_XI13/Mm1_s
+ N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=3.5e-07 AD=2.629e-13 AS=2.629e-13
+ PD=1.77e-06 PS=1.77e-06
mXI25/XI1/MM8 N_LFSR8_XI25/XI1/MM8_d N_LFSR8_BAR_XI25/XI1/MM8_g
+ N_VDD_XI25/XI1/MM8_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI18/XI1/MM4 N_XI18/XI1/NET8_XI18/XI1/MM4_d N_CLK_XI18/XI1/MM4_g
+ N_XI18/XI1/NET39_XI18/XI1/MM4_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07
+ AD=3.43e-13 AS=8.75e-14 PD=1.68e-06 PS=2.5e-07
mXI18/XI4/MM4 N_XI18/XI4/NET8_XI18/XI4/MM4_d N_CLK_XI18/XI4/MM4_g
+ N_XI18/XI4/NET39_XI18/XI4/MM4_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07
+ W=7e-07 AD=3.43e-13 AS=8.75e-14 PD=1.68e-06 PS=2.5e-07
mXI18/XI1/MM5 N_XI18/XI1/NET39_XI18/XI1/MM5_d N_XI18/PREBIT0_XI18/XI1/MM5_g
+ N_VDD_XI18/XI1/MM5_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=8.75e-14
+ AS=3.43e-13 PD=2.5e-07 PS=1.68e-06
mXI18/XI4/MM5 N_XI18/XI4/NET39_XI18/XI4/MM5_d N_XI18/PREBIT1_XI18/XI4/MM5_g
+ N_VDD_XI18/XI4/MM5_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07 W=7e-07
+ AD=8.75e-14 AS=3.43e-13 PD=2.5e-07 PS=1.68e-06
mXI25/XI6/MM7 N_LFSR2_BAR_XI25/XI6/MM7_d N_XI25/XI6/NET31_XI25/XI6/MM7_g
+ N_VDD_XI25/XI6/MM7_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=7e-07 AD=7.07e-13
+ AS=3.43e-13 PD=2.72e-06 PS=1.68e-06
mXI25/XI1/MM7 N_LFSR8_BAR_XI25/XI1/MM7_d N_XI25/XI1/NET22_XI25/XI1/MM7_g
+ N_VDD_XI25/XI1/MM7_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI17/XI7/MM8 N_XI17/A0_XI17/XI7/MM8_d N_XI17/A0BAR_XI17/XI7/MM8_g
+ N_VDD_XI17/XI7/MM8_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI17/XI6/MM8 N_XI17/A1_XI17/XI6/MM8_d N_XI17/A1BAR_XI17/XI6/MM8_g
+ N_VDD_XI17/XI6/MM8_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI25/XI6/MM8 N_LFSR2_XI25/XI6/MM8_d N_LFSR2_BAR_XI25/XI6/MM8_g
+ N_VDD_XI25/XI6/MM8_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI25/XI1/MM6 N_XI25/XI1/NET22_XI25/XI1/MM6_d N_CLK_XI25/XI1/MM6_g
+ N_VDD_XI25/XI1/MM6_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI17/XI7/MM11 N_XI17/A0BAR_XI17/XI7/MM11_d N_RSTOBAR_XI17/XI7/MM11_g
+ N_VDD_XI17/XI7/MM11_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI17/XI6/MM11 N_XI17/A1BAR_XI17/XI6/MM11_d N_RSTOBAR_XI17/XI6/MM11_g
+ N_VDD_XI17/XI6/MM11_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI18/XI6/MM8 N_XI18/PREBIT0_XI18/XI6/MM8_d N_XI18/NET40_XI18/XI6/MM8_g
+ N_VDD_XI18/XI6/MM8_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI18/XI9/MM8 N_XI18/PREBIT1_XI18/XI9/MM8_d N_XI18/NET47_XI18/XI9/MM8_g
+ N_VDD_XI18/XI9/MM8_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07 W=7e-07
+ AD=3.43e-13 AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI25/XI1/MM4 N_XI25/XI1/NET6_XI25/XI1/MM4_d N_CLK_XI25/XI1/MM4_g
+ N_XI25/XI1/NET33_XI25/XI1/MM4_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=2.25e-13 PD=2.78e-06 PS=2.5e-07
mXI17/XI7/MM7 N_XI17/A0BAR_XI17/XI7/MM7_d N_XI17/XI7/NET24_XI17/XI7/MM7_g
+ N_VDD_XI17/XI7/MM7_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=6.44e-13
+ AS=3.43e-13 PD=2.54e-06 PS=1.68e-06
mXI17/XI6/MM7 N_XI17/A1BAR_XI17/XI6/MM7_d N_XI17/XI6/NET24_XI17/XI6/MM7_g
+ N_VDD_XI17/XI6/MM7_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=7e-07 AD=6.44e-13
+ AS=3.43e-13 PD=2.54e-06 PS=1.68e-06
mXI25/XI1/MM5 N_XI25/XI1/NET33_XI25/XI1/MM5_d N_LFSR7_XI25/XI1/MM5_g
+ N_VDD_XI25/XI1/MM5_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=2.25e-13
+ AS=8.82e-13 PD=2.5e-07 PS=2.78e-06
mXI18/XI6/MM7 N_XI18/NET40_XI18/XI6/MM7_d N_XI18/XI6/NET31_XI18/XI6/MM7_g
+ N_VDD_XI18/XI6/MM7_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=7.07e-13
+ AS=3.43e-13 PD=2.72e-06 PS=1.68e-06
mXI18/XI9/MM7 N_XI18/NET47_XI18/XI9/MM7_d N_XI18/XI9/NET31_XI18/XI9/MM7_g
+ N_VDD_XI18/XI9/MM7_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07 W=7e-07
+ AD=7.07e-13 AS=3.43e-13 PD=2.72e-06 PS=1.68e-06
mXI25/XI3/MM8 N_LFSR7_XI25/XI3/MM8_d N_LFSR7_BAR_XI25/XI3/MM8_g
+ N_VDD_XI25/XI3/MM8_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI17/XI7/MM6 N_XI17/XI7/NET24_XI17/XI7/MM6_d N_CLK_XI17/XI7/MM6_g
+ N_VDD_XI17/XI7/MM6_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI17/XI6/MM6 N_XI17/XI6/NET24_XI17/XI6/MM6_d N_CLK_XI17/XI6/MM6_g
+ N_VDD_XI17/XI6/MM6_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=3.43e-13 PD=1.68e-06 PS=1.68e-06
mXI25/XI18/MM5 N_XI25/XI18/NET33_XI25/XI18/MM5_d N_LFSR2_XI25/XI18/MM5_g
+ N_VDD_XI25/XI18/MM5_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06
+ AD=2.25e-13 AS=8.82e-13 PD=2.5e-07 PS=2.78e-06
mXI25/XI18/MM4 N_XI25/XI18/NET6_XI25/XI18/MM4_d N_CLK_XI25/XI18/MM4_g
+ N_XI25/XI18/NET33_XI25/XI18/MM4_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07
+ W=1.8e-06 AD=8.82e-13 AS=2.25e-13 PD=2.78e-06 PS=2.5e-07
mXI25/XI3/MM7 N_LFSR7_BAR_XI25/XI3/MM7_d N_XI25/XI3/NET22_XI25/XI3/MM7_g
+ N_VDD_XI25/XI3/MM7_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI17/XI7/MM4 N_XI17/XI7/NET8_XI17/XI7/MM4_d N_CLK_XI17/XI7/MM4_g
+ N_XI17/XI7/NET39_XI17/XI7/MM4_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07
+ AD=3.43e-13 AS=8.75e-14 PD=1.68e-06 PS=2.5e-07
mXI17/XI6/MM4 N_XI17/XI6/NET8_XI17/XI6/MM4_d N_CLK_XI17/XI6/MM4_g
+ N_XI17/XI6/NET39_XI17/XI6/MM4_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=7e-07
+ AD=3.43e-13 AS=8.75e-14 PD=1.68e-06 PS=2.5e-07
mXI18/XI6/MM6 N_XI18/XI6/NET31_XI18/XI6/MM6_d N_CLK_XI18/XI6/MM6_g
+ N_VDD_XI18/XI6/MM6_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=3.43e-13
+ AS=4.935e-13 PD=1.68e-06 PS=2.11e-06
mXI18/XI9/MM6 N_XI18/XI9/NET31_XI18/XI9/MM6_d N_CLK_XI18/XI9/MM6_g
+ N_VDD_XI18/XI9/MM6_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07 W=7e-07
+ AD=3.43e-13 AS=4.935e-13 PD=1.68e-06 PS=2.11e-06
mXI17/XI7/MM5 N_XI17/XI7/NET39_XI17/XI7/MM5_d N_NET083_XI17/XI7/MM5_g
+ N_VDD_XI17/XI7/MM5_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=8.75e-14
+ AS=3.43e-13 PD=2.5e-07 PS=1.68e-06
mXI17/XI6/MM5 N_XI17/XI6/NET39_XI17/XI6/MM5_d N_NET082_XI17/XI6/MM5_g
+ N_VDD_XI17/XI6/MM5_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=7e-07 AD=8.75e-14
+ AS=3.43e-13 PD=2.5e-07 PS=1.68e-06
mXI25/XI18/MM6 N_XI25/XI18/NET22_XI25/XI18/MM6_d N_CLK_XI25/XI18/MM6_g
+ N_VDD_XI25/XI18/MM6_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI3/MM6 N_XI25/XI3/NET22_XI25/XI3/MM6_d N_CLK_XI25/XI3/MM6_g
+ N_VDD_XI25/XI3/MM6_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=8.82e-13
+ AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI18/XI6/MM4 N_XI18/XI6/NET47_XI18/XI6/MM4_d N_CLK_XI18/XI6/MM4_g
+ N_XI18/XI6/NET26_XI18/XI6/MM4_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07
+ AD=4.095e-13 AS=8.75e-14 PD=1.87e-06 PS=2.5e-07
mXI18/XI9/MM4 N_XI18/XI9/NET47_XI18/XI9/MM4_d N_CLK_XI18/XI9/MM4_g
+ N_XI18/XI9/NET26_XI18/XI9/MM4_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07
+ W=7e-07 AD=4.095e-13 AS=8.75e-14 PD=1.87e-06 PS=2.5e-07
mXI17/XI1/XI2/MM1 N_XI17/NET13_XI17/XI1/XI2/MM1_d N_LFSR7_XI17/XI1/XI2/MM1_g
+ N_NET082_XI17/XI1/XI2/MM1_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI4/XI2/MM1 N_XI17/NET024_XI17/XI4/XI2/MM1_d
+ N_LFSR7_BAR_XI17/XI4/XI2/MM1_g N_NET083_XI17/XI4/XI2/MM1_s
+ N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI18/XI6/MM5 N_XI18/XI6/NET26_XI18/XI6/MM5_d N_NET071_XI18/XI6/MM5_g
+ N_VDD_XI18/XI6/MM5_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=7e-07 AD=8.75e-14
+ AS=3.43e-13 PD=2.5e-07 PS=1.68e-06
mXI18/XI9/MM5 N_XI18/XI9/NET26_XI18/XI9/MM5_d N_NET070_XI18/XI9/MM5_g
+ N_VDD_XI18/XI9/MM5_s N_VDD_XI18/XI3/XI1/MM1_b P_18 L=1.8e-07 W=7e-07
+ AD=8.75e-14 AS=3.43e-13 PD=2.5e-07 PS=1.68e-06
mXI25/XI18/MM7 N_LFSR3_BAR_XI25/XI18/MM7_d N_XI25/XI18/NET22_XI25/XI18/MM7_g
+ N_VDD_XI25/XI18/MM7_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI3/MM4 N_XI25/XI3/NET6_XI25/XI3/MM4_d N_CLK_XI25/XI3/MM4_g
+ N_XI25/XI3/NET33_XI25/XI3/MM4_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=2.25e-13 PD=2.78e-06 PS=2.5e-07
mXI17/XI1/XI1/MM1 N_XI17/A1BAR_XI17/XI1/XI1/MM1_d N_LFSR7_BAR_XI17/XI1/XI1/MM1_g
+ N_NET082_XI17/XI1/XI1/MM1_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI4/XI1/MM1 N_XI17/A0BAR_XI17/XI4/XI1/MM1_d N_LFSR7_XI17/XI4/XI1/MM1_g
+ N_NET083_XI17/XI4/XI1/MM1_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI3/MM5 N_XI25/XI3/NET33_XI25/XI3/MM5_d N_LFSR6_XI25/XI3/MM5_g
+ N_VDD_XI25/XI3/MM5_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06 AD=2.25e-13
+ AS=8.82e-13 PD=2.5e-07 PS=2.78e-06
mXI25/XI18/MM8 N_LFSR3_XI25/XI18/MM8_d N_LFSR3_BAR_XI25/XI18/MM8_g
+ N_VDD_XI25/XI18/MM8_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI14/MM8 N_LFSR6_XI25/XI14/MM8_d N_LFSR6_BAR_XI25/XI14/MM8_g
+ N_VDD_XI25/XI14/MM8_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI2/XI3/MM1 N_LFSR3_XI25/XI2/XI3/MM1_d N_LFSR10_XI25/XI2/XI3/MM1_g
+ N_XI25/NET62_XI25/XI2/XI3/MM1_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI2/XI2/MM1 N_XI17/A1_XI17/XI2/XI2/MM1_d N_LFSR5_XI17/XI2/XI2/MM1_g
+ N_XI17/NET13_XI17/XI2/XI2/MM1_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI3/XI2/MM1 N_XI17/A0_XI17/XI3/XI2/MM1_d N_LFSR5_XI17/XI3/XI2/MM1_g
+ N_XI17/NET024_XI17/XI3/XI2/MM1_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI14/MM7 N_LFSR6_BAR_XI25/XI14/MM7_d N_XI25/XI14/NET22_XI25/XI14/MM7_g
+ N_VDD_XI25/XI14/MM7_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI5/XI0/XI0/XI2/MM1 N_NET071_XI5/XI0/XI0/XI2/MM1_d N_M0_XI5/XI0/XI0/XI2/MM1_g
+ N_XI5/XI0/NET40_XI5/XI0/XI0/XI2/MM1_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI0/XI1/MM1 N_NET089_XI5/XI0/XI0/XI1/MM1_d
+ N_M0_BAR_XI5/XI0/XI0/XI1/MM1_g N_XI5/XI0/NET40_XI5/XI0/XI0/XI1/MM1_s
+ N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI7/XI1/MM1 N_NET087_XI5/XI0/XI7/XI1/MM1_d
+ N_M0_BAR_XI5/XI0/XI7/XI1/MM1_g N_XI5/XI0/NET33_XI5/XI0/XI7/XI1/MM1_s
+ N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI7/XI2/MM1 N_NET070_XI5/XI0/XI7/XI2/MM1_d N_M0_XI5/XI0/XI7/XI2/MM1_g
+ N_XI5/XI0/NET33_XI5/XI0/XI7/XI2/MM1_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07
+ W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI2/XI2/MM1 N_LFSR3_BAR_XI25/XI2/XI2/MM1_d N_LFSR10_BAR_XI25/XI2/XI2/MM1_g
+ N_XI25/NET62_XI25/XI2/XI2/MM1_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI2/XI1/MM1 N_LFSR6_XI17/XI2/XI1/MM1_d N_LFSR5_BAR_XI17/XI2/XI1/MM1_g
+ N_XI17/NET13_XI17/XI2/XI1/MM1_s N_VDD_XI4/XI8/MM5_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI17/XI3/XI1/MM1 N_LFSR6_XI17/XI3/XI1/MM1_d N_LFSR5_BAR_XI17/XI3/XI1/MM1_g
+ N_XI17/NET024_XI17/XI3/XI1/MM1_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI14/MM6 N_XI25/XI14/NET22_XI25/XI14/MM6_d N_CLK_XI25/XI14/MM6_g
+ N_VDD_XI25/XI14/MM6_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI16/MM5 N_XI25/XI16/NET33_XI25/XI16/MM5_d N_XI25/NET62_XI25/XI16/MM5_g
+ N_VDD_XI25/XI16/MM5_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06
+ AD=2.25e-13 AS=8.82e-13 PD=2.5e-07 PS=2.78e-06
mXI25/XI16/MM4 N_XI25/XI16/NET6_XI25/XI16/MM4_d N_CLK_XI25/XI16/MM4_g
+ N_XI25/XI16/NET33_XI25/XI16/MM4_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07
+ W=1.8e-06 AD=8.82e-13 AS=2.25e-13 PD=2.78e-06 PS=2.5e-07
mXI25/XI14/MM4 N_XI25/XI14/NET6_XI25/XI14/MM4_d N_CLK_XI25/XI14/MM4_g
+ N_XI25/XI14/NET33_XI25/XI14/MM4_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07
+ W=1.8e-06 AD=8.82e-13 AS=2.25e-13 PD=2.78e-06 PS=2.5e-07
mXI25/XI14/MM5 N_XI25/XI14/NET33_XI25/XI14/MM5_d N_LFSR5_XI25/XI14/MM5_g
+ N_VDD_XI25/XI14/MM5_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06
+ AD=2.25e-13 AS=8.82e-13 PD=2.5e-07 PS=2.78e-06
mXI25/XI16/MM6 N_XI25/XI16/NET22_XI25/XI16/MM6_d N_CLK_XI25/XI16/MM6_g
+ N_VDD_XI25/XI16/MM6_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI5/XI0/XI2/XI2/MM1 N_XI5/XI0/NET54_XI5/XI0/XI2/XI2/MM1_d
+ N_M1_XI5/XI0/XI2/XI2/MM1_g N_XI5/NET64_XI5/XI0/XI2/XI2/MM1_s
+ N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI2/XI1/MM1 N_XI5/XI0/NET40_XI5/XI0/XI2/XI1/MM1_d
+ N_M1_BAR_XI5/XI0/XI2/XI1/MM1_g N_XI5/NET64_XI5/XI0/XI2/XI1/MM1_s
+ N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI8/XI1/MM1 N_XI5/XI0/NET33_XI5/XI0/XI8/XI1/MM1_d
+ N_M1_BAR_XI5/XI0/XI8/XI1/MM1_g N_XI5/NET63_XI5/XI0/XI8/XI1/MM1_s
+ N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI8/XI2/MM1 N_XI5/XI0/NET19_XI5/XI0/XI8/XI2/MM1_d
+ N_M1_XI5/XI0/XI8/XI2/MM1_g N_XI5/NET63_XI5/XI0/XI8/XI2/MM1_s
+ N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI25/XI15/MM8 N_LFSR5_XI25/XI15/MM8_d N_LFSR5_BAR_XI25/XI15/MM8_g
+ N_VDD_XI25/XI15/MM8_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI16/MM7 N_LFSR4_BAR_XI25/XI16/MM7_d N_XI25/XI16/NET22_XI25/XI16/MM7_g
+ N_VDD_XI25/XI16/MM7_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI5/XI0/XI9/XI2/MM1 N_LFSR8_XI5/XI0/XI9/XI2/MM1_d N_M0_XI5/XI0/XI9/XI2/MM1_g
+ N_XI5/XI0/NET19_XI5/XI0/XI9/XI2/MM1_s N_VDD_XI5/XI0/XI9/XI2/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI9/XI1/MM1 N_NET082_XI5/XI0/XI9/XI1/MM1_d
+ N_M0_BAR_XI5/XI0/XI9/XI1/MM1_g N_XI5/XI0/NET19_XI5/XI0/XI9/XI1/MM1_s
+ N_VDD_XI5/XI0/XI9/XI2/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI1/XI1/MM1 N_NET083_XI5/XI0/XI1/XI1/MM1_d
+ N_M0_BAR_XI5/XI0/XI1/XI1/MM1_g N_XI5/XI0/NET54_XI5/XI0/XI1/XI1/MM1_s
+ N_VDD_XI5/XI0/XI9/XI2/MM1_b P_18 L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13
+ PD=1.48e-06 PS=1.48e-06
mXI5/XI0/XI1/XI2/MM1 N_LFSR3_XI5/XI0/XI1/XI2/MM1_d N_M0_XI5/XI0/XI1/XI2/MM1_g
+ N_XI5/XI0/NET54_XI5/XI0/XI1/XI2/MM1_s N_VDD_XI5/XI0/XI9/XI2/MM1_b P_18
+ L=1.8e-07 W=5e-07 AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
mXI25/XI15/MM7 N_LFSR5_BAR_XI25/XI15/MM7_d N_XI25/XI15/NET22_XI25/XI15/MM7_g
+ N_VDD_XI25/XI15/MM7_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI25/XI16/MM8 N_LFSR4_XI25/XI16/MM8_d N_LFSR4_BAR_XI25/XI16/MM8_g
+ N_VDD_XI25/XI16/MM8_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI5/XI2/Mm1 N_XI5/NET42_XI5/XI2/Mm1_d N_XI5/NET64_XI5/XI2/Mm1_g
+ N_VDD_XI5/XI2/Mm1_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=3.5e-07 AD=2.629e-13
+ AS=2.629e-13 PD=1.77e-06 PS=1.77e-06
mXI5/XI3/Mm1 N_XI5/NET38_XI5/XI3/Mm1_d N_XI5/NET63_XI5/XI3/Mm1_g
+ N_VDD_XI5/XI3/Mm1_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=3.5e-07 AD=2.629e-13
+ AS=2.629e-13 PD=1.77e-06 PS=1.77e-06
mXI25/XI15/MM6 N_XI25/XI15/NET22_XI25/XI15/MM6_d N_CLK_XI25/XI15/MM6_g
+ N_VDD_XI25/XI15/MM6_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06
+ AD=8.82e-13 AS=8.82e-13 PD=2.78e-06 PS=2.78e-06
mXI7/Mm1 N_M0_BAR_XI7/Mm1_d N_M0_XI7/Mm1_g N_VDD_XI7/Mm1_s
+ N_VDD_XI5/XI0/XI9/XI2/MM1_b P_18 L=1.8e-07 W=3.5e-07 AD=2.629e-13 AS=2.629e-13
+ PD=1.77e-06 PS=1.77e-06
mXI8/Mm1 N_M1_BAR_XI8/Mm1_d N_M1_XI8/Mm1_g N_VDD_XI8/Mm1_s
+ N_VDD_XI5/XI0/XI9/XI2/MM1_b P_18 L=1.8e-07 W=3.5e-07 AD=2.629e-13 AS=2.629e-13
+ PD=1.77e-06 PS=1.77e-06
mXI5/XI1/MM13 N_VDD_XI5/XI1/MM13_d N_XI5/NET42_XI5/XI1/MM13_g
+ N_XI5/XI1/NET72_XI5/XI1/MM13_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=2.5e-07
+ AD=2.509e-13 AS=3.5e-14 PD=1.87e-06 PS=2.8e-07
mXI5/XI1/MM8 N_VDD_XI5/XI1/MM8_d N_XI5/NET64_XI5/XI1/MM8_g
+ N_XI5/XI1/NET60_XI5/XI1/MM8_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=2.5e-07
+ AD=2.509e-13 AS=3.5e-14 PD=1.87e-06 PS=2.8e-07
mXI5/XI1/MM2 N_VDD_XI5/XI1/MM2_d N_XI5/NET64_XI5/XI1/MM2_g
+ N_XI5/XI1/NET44_XI5/XI1/MM2_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=2.5e-07
+ AD=2.509e-13 AS=3.5e-14 PD=1.87e-06 PS=2.8e-07
mXI5/XI1/MM5 N_VDD_XI5/XI1/MM5_d N_XI5/NET42_XI5/XI1/MM5_g
+ N_XI5/XI1/NET56_XI5/XI1/MM5_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=2.5e-07
+ AD=2.509e-13 AS=3.5e-14 PD=1.87e-06 PS=2.8e-07
mXI5/XI1/MM12 N_XI5/XI1/NET72_XI5/XI1/MM12_d N_XI5/NET38_XI5/XI1/MM12_g
+ N_CH3_XI5/XI1/MM12_s N_VDD_XI25/XI4/MM8_b P_18 L=1.8e-07 W=2.5e-07 AD=3.5e-14
+ AS=2.509e-13 PD=2.8e-07 PS=1.87e-06
mXI5/XI1/MM9 N_XI5/XI1/NET60_XI5/XI1/MM9_d N_XI5/NET38_XI5/XI1/MM9_g
+ N_CH2_XI5/XI1/MM9_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=2.5e-07 AD=3.5e-14
+ AS=2.509e-13 PD=2.8e-07 PS=1.87e-06
mXI5/XI1/MM3 N_XI5/XI1/NET44_XI5/XI1/MM3_d N_XI5/NET63_XI5/XI1/MM3_g
+ N_CH0_XI5/XI1/MM3_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=2.5e-07 AD=3.5e-14
+ AS=2.509e-13 PD=2.8e-07 PS=1.87e-06
mXI5/XI1/MM4 N_XI5/XI1/NET56_XI5/XI1/MM4_d N_XI5/NET63_XI5/XI1/MM4_g
+ N_CH1_XI5/XI1/MM4_s N_VDD_XI4/XI10/MM8_b P_18 L=1.8e-07 W=2.5e-07 AD=3.5e-14
+ AS=2.509e-13 PD=2.8e-07 PS=1.87e-06
mXI25/XI15/MM4 N_XI25/XI15/NET6_XI25/XI15/MM4_d N_CLK_XI25/XI15/MM4_g
+ N_XI25/XI15/NET33_XI25/XI15/MM4_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07
+ W=1.8e-06 AD=8.82e-13 AS=2.25e-13 PD=2.78e-06 PS=2.5e-07
mXI25/XI15/MM5 N_XI25/XI15/NET33_XI25/XI15/MM5_d N_LFSR4_XI25/XI15/MM5_g
+ N_VDD_XI25/XI15/MM5_s N_VDD_XI25/XI4/MM7_b P_18 L=1.8e-07 W=1.8e-06
+ AD=2.25e-13 AS=8.82e-13 PD=2.5e-07 PS=2.78e-06
*
.include "RIS.pex.spi.RIS.pxi"
*
.ends
*
*
